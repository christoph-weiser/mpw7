.subckt user_analog_project_wrapper vdda1 vdda2 vssa1 vssa2 vccd1 vccd2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_stb_i wbs_cyc_i wbs_we_i wbs_sel_i[3] wbs_sel_i[2] wbs_sel_i[1] wbs_sel_i[0] wbs_dat_i[31]
+ wbs_dat_i[30] wbs_dat_i[29] wbs_dat_i[28] wbs_dat_i[27] wbs_dat_i[26] wbs_dat_i[25] wbs_dat_i[24] wbs_dat_i[23]
+ wbs_dat_i[22] wbs_dat_i[21] wbs_dat_i[20] wbs_dat_i[19] wbs_dat_i[18] wbs_dat_i[17] wbs_dat_i[16] wbs_dat_i[15]
+ wbs_dat_i[14] wbs_dat_i[13] wbs_dat_i[12] wbs_dat_i[11] wbs_dat_i[10] wbs_dat_i[9] wbs_dat_i[8] wbs_dat_i[7]
+ wbs_dat_i[6] wbs_dat_i[5] wbs_dat_i[4] wbs_dat_i[3] wbs_dat_i[2] wbs_dat_i[1] wbs_dat_i[0] wbs_adr_i[31]
+ wbs_adr_i[30] wbs_adr_i[29] wbs_adr_i[28] wbs_adr_i[27] wbs_adr_i[26] wbs_adr_i[25] wbs_adr_i[24] wbs_adr_i[23]
+ wbs_adr_i[22] wbs_adr_i[21] wbs_adr_i[20] wbs_adr_i[19] wbs_adr_i[18] wbs_adr_i[17] wbs_adr_i[16] wbs_adr_i[15]
+ wbs_adr_i[14] wbs_adr_i[13] wbs_adr_i[12] wbs_adr_i[11] wbs_adr_i[10] wbs_adr_i[9] wbs_adr_i[8] wbs_adr_i[7]
+ wbs_adr_i[6] wbs_adr_i[5] wbs_adr_i[4] wbs_adr_i[3] wbs_adr_i[2] wbs_adr_i[1] wbs_adr_i[0] wbs_ack_o
+ wbs_dat_o[31] wbs_dat_o[30] wbs_dat_o[29] wbs_dat_o[28] wbs_dat_o[27] wbs_dat_o[26] wbs_dat_o[25] wbs_dat_o[24]
+ wbs_dat_o[23] wbs_dat_o[22] wbs_dat_o[21] wbs_dat_o[20] wbs_dat_o[19] wbs_dat_o[18] wbs_dat_o[17] wbs_dat_o[16]
+ wbs_dat_o[15] wbs_dat_o[14] wbs_dat_o[13] wbs_dat_o[12] wbs_dat_o[11] wbs_dat_o[10] wbs_dat_o[9] wbs_dat_o[8]
+ wbs_dat_o[7] wbs_dat_o[6] wbs_dat_o[5] wbs_dat_o[4] wbs_dat_o[3] wbs_dat_o[2] wbs_dat_o[1] wbs_dat_o[0]
+ la_data_in[127] la_data_in[126] la_data_in[125] la_data_in[124] la_data_in[123] la_data_in[122] la_data_in[121]
+ la_data_in[120] la_data_in[119] la_data_in[118] la_data_in[117] la_data_in[116] la_data_in[115] la_data_in[114]
+ la_data_in[113] la_data_in[112] la_data_in[111] la_data_in[110] la_data_in[109] la_data_in[108] la_data_in[107]
+ la_data_in[106] la_data_in[105] la_data_in[104] la_data_in[103] la_data_in[102] la_data_in[101] la_data_in[100]
+ la_data_in[99] la_data_in[98] la_data_in[97] la_data_in[96] la_data_in[95] la_data_in[94] la_data_in[93]
+ la_data_in[92] la_data_in[91] la_data_in[90] la_data_in[89] la_data_in[88] la_data_in[87] la_data_in[86]
+ la_data_in[85] la_data_in[84] la_data_in[83] la_data_in[82] la_data_in[81] la_data_in[80] la_data_in[79]
+ la_data_in[78] la_data_in[77] la_data_in[76] la_data_in[75] la_data_in[74] la_data_in[73] la_data_in[72]
+ la_data_in[71] la_data_in[70] la_data_in[69] la_data_in[68] la_data_in[67] la_data_in[66] la_data_in[65]
+ la_data_in[64] la_data_in[63] la_data_in[62] la_data_in[61] la_data_in[60] la_data_in[59] la_data_in[58]
+ la_data_in[57] la_data_in[56] la_data_in[55] la_data_in[54] la_data_in[53] la_data_in[52] la_data_in[51]
+ la_data_in[50] la_data_in[49] la_data_in[48] la_data_in[47] la_data_in[46] la_data_in[45] la_data_in[44]
+ la_data_in[43] la_data_in[42] la_data_in[41] la_data_in[40] la_data_in[39] la_data_in[38] la_data_in[37]
+ la_data_in[36] la_data_in[35] la_data_in[34] la_data_in[33] la_data_in[32] la_data_in[31] la_data_in[30]
+ la_data_in[29] la_data_in[28] la_data_in[27] la_data_in[26] la_data_in[25] la_data_in[24] la_data_in[23]
+ la_data_in[22] la_data_in[21] la_data_in[20] la_data_in[19] la_data_in[18] la_data_in[17] la_data_in[16]
+ la_data_in[15] la_data_in[14] la_data_in[13] la_data_in[12] la_data_in[11] la_data_in[10] la_data_in[9]
+ la_data_in[8] la_data_in[7] la_data_in[6] la_data_in[5] la_data_in[4] la_data_in[3] la_data_in[2] la_data_in[1]
+ la_data_in[0] la_data_out[127] la_data_out[126] la_data_out[125] la_data_out[124] la_data_out[123]
+ la_data_out[122] la_data_out[121] la_data_out[120] la_data_out[119] la_data_out[118] la_data_out[117]
+ la_data_out[116] la_data_out[115] la_data_out[114] la_data_out[113] la_data_out[112] la_data_out[111]
+ la_data_out[110] la_data_out[109] la_data_out[108] la_data_out[107] la_data_out[106] la_data_out[105]
+ la_data_out[104] la_data_out[103] la_data_out[102] la_data_out[101] la_data_out[100] la_data_out[99] la_data_out[98]
+ la_data_out[97] la_data_out[96] la_data_out[95] la_data_out[94] la_data_out[93] la_data_out[92] la_data_out[91]
+ la_data_out[90] la_data_out[89] la_data_out[88] la_data_out[87] la_data_out[86] la_data_out[85] la_data_out[84]
+ la_data_out[83] la_data_out[82] la_data_out[81] la_data_out[80] la_data_out[79] la_data_out[78] la_data_out[77]
+ la_data_out[76] la_data_out[75] la_data_out[74] la_data_out[73] la_data_out[72] la_data_out[71] la_data_out[70]
+ la_data_out[69] la_data_out[68] la_data_out[67] la_data_out[66] la_data_out[65] la_data_out[64] la_data_out[63]
+ la_data_out[62] la_data_out[61] la_data_out[60] la_data_out[59] la_data_out[58] la_data_out[57] la_data_out[56]
+ la_data_out[55] la_data_out[54] la_data_out[53] la_data_out[52] la_data_out[51] la_data_out[50] la_data_out[49]
+ la_data_out[48] la_data_out[47] la_data_out[46] la_data_out[45] la_data_out[44] la_data_out[43] la_data_out[42]
+ la_data_out[41] la_data_out[40] la_data_out[39] la_data_out[38] la_data_out[37] la_data_out[36] la_data_out[35]
+ la_data_out[34] la_data_out[33] la_data_out[32] la_data_out[31] la_data_out[30] la_data_out[29] la_data_out[28]
+ la_data_out[27] la_data_out[26] la_data_out[25] la_data_out[24] la_data_out[23] la_data_out[22] la_data_out[21]
+ la_data_out[20] la_data_out[19] la_data_out[18] la_data_out[17] la_data_out[16] la_data_out[15] la_data_out[14]
+ la_data_out[13] la_data_out[12] la_data_out[11] la_data_out[10] la_data_out[9] la_data_out[8] la_data_out[7]
+ la_data_out[6] la_data_out[5] la_data_out[4] la_data_out[3] la_data_out[2] la_data_out[1] la_data_out[0] io_in[26]
+ io_in[25] io_in[24] io_in[23] io_in[22] io_in[21] io_in[20] io_in[19] io_in[18] io_in[17] io_in[16] io_in[15]
+ io_in[14] io_in[13] io_in[12] io_in[11] io_in[10] io_in[9] io_in[8] io_in[7] io_in[6] io_in[5] io_in[4]
+ io_in[3] io_in[2] io_in[1] io_in[0] io_in_3v3[26] io_in_3v3[25] io_in_3v3[24] io_in_3v3[23] io_in_3v3[22]
+ io_in_3v3[21] io_in_3v3[20] io_in_3v3[19] io_in_3v3[18] io_in_3v3[17] io_in_3v3[16] io_in_3v3[15] io_in_3v3[14]
+ io_in_3v3[13] io_in_3v3[12] io_in_3v3[11] io_in_3v3[10] io_in_3v3[9] io_in_3v3[8] io_in_3v3[7] io_in_3v3[6]
+ io_in_3v3[5] io_in_3v3[4] io_in_3v3[3] io_in_3v3[2] io_in_3v3[1] io_in_3v3[0] user_clock2 io_out[26] io_out[25]
+ io_out[24] io_out[23] io_out[22] io_out[21] io_out[20] io_out[19] io_out[18] io_out[17] io_out[16] io_out[15]
+ io_out[14] io_out[13] io_out[12] io_out[11] io_out[10] io_out[9] io_out[8] io_out[7] io_out[6] io_out[5]
+ io_out[4] io_out[3] io_out[2] io_out[1] io_out[0] io_oeb[26] io_oeb[25] io_oeb[24] io_oeb[23] io_oeb[22]
+ io_oeb[21] io_oeb[20] io_oeb[19] io_oeb[18] io_oeb[17] io_oeb[16] io_oeb[15] io_oeb[14] io_oeb[13] io_oeb[12]
+ io_oeb[11] io_oeb[10] io_oeb[9] io_oeb[8] io_oeb[7] io_oeb[6] io_oeb[5] io_oeb[4] io_oeb[3] io_oeb[2]
+ io_oeb[1] io_oeb[0] gpio_analog[17] gpio_analog[16] gpio_analog[15] gpio_analog[14] gpio_analog[13]
+ gpio_analog[12] gpio_analog[11] gpio_analog[10] gpio_analog[9] gpio_analog[8] gpio_analog[7] gpio_analog[6]
+ gpio_analog[5] gpio_analog[4] gpio_analog[3] gpio_analog[2] gpio_analog[1] gpio_analog[0] gpio_noesd[17]
+ gpio_noesd[16] gpio_noesd[15] gpio_noesd[14] gpio_noesd[13] gpio_noesd[12] gpio_noesd[11] gpio_noesd[10]
+ gpio_noesd[9] gpio_noesd[8] gpio_noesd[7] gpio_noesd[6] gpio_noesd[5] gpio_noesd[4] gpio_noesd[3] gpio_noesd[2]
+ gpio_noesd[1] gpio_noesd[0] io_analog[10] io_analog[9] io_analog[8] io_analog[7] io_analog[6] io_analog[5]
+ io_analog[4] io_analog[3] io_analog[2] io_analog[1] io_analog[0] io_clamp_high[2] io_clamp_high[1]
+ io_clamp_high[0] io_clamp_low[2] io_clamp_low[1] io_clamp_low[0] user_irq[2] user_irq[1] user_irq[0] la_oenb[127]
+ la_oenb[126] la_oenb[125] la_oenb[124] la_oenb[123] la_oenb[122] la_oenb[121] la_oenb[120] la_oenb[119]
+ la_oenb[118] la_oenb[117] la_oenb[116] la_oenb[115] la_oenb[114] la_oenb[113] la_oenb[112] la_oenb[111]
+ la_oenb[110] la_oenb[109] la_oenb[108] la_oenb[107] la_oenb[106] la_oenb[105] la_oenb[104] la_oenb[103]
+ la_oenb[102] la_oenb[101] la_oenb[100] la_oenb[99] la_oenb[98] la_oenb[97] la_oenb[96] la_oenb[95] la_oenb[94]
+ la_oenb[93] la_oenb[92] la_oenb[91] la_oenb[90] la_oenb[89] la_oenb[88] la_oenb[87] la_oenb[86] la_oenb[85]
+ la_oenb[84] la_oenb[83] la_oenb[82] la_oenb[81] la_oenb[80] la_oenb[79] la_oenb[78] la_oenb[77] la_oenb[76]
+ la_oenb[75] la_oenb[74] la_oenb[73] la_oenb[72] la_oenb[71] la_oenb[70] la_oenb[69] la_oenb[68] la_oenb[67]
+ la_oenb[66] la_oenb[65] la_oenb[64] la_oenb[63] la_oenb[62] la_oenb[61] la_oenb[60] la_oenb[59] la_oenb[58]
+ la_oenb[57] la_oenb[56] la_oenb[55] la_oenb[54] la_oenb[53] la_oenb[52] la_oenb[51] la_oenb[50] la_oenb[49]
+ la_oenb[48] la_oenb[47] la_oenb[46] la_oenb[45] la_oenb[44] la_oenb[43] la_oenb[42] la_oenb[41] la_oenb[40]
+ la_oenb[39] la_oenb[38] la_oenb[37] la_oenb[36] la_oenb[35] la_oenb[34] la_oenb[33] la_oenb[32] la_oenb[31]
+ la_oenb[30] la_oenb[29] la_oenb[28] la_oenb[27] la_oenb[26] la_oenb[25] la_oenb[24] la_oenb[23] la_oenb[22]
+ la_oenb[21] la_oenb[20] la_oenb[19] la_oenb[18] la_oenb[17] la_oenb[16] la_oenb[15] la_oenb[14] la_oenb[13]
+ la_oenb[12] la_oenb[11] la_oenb[10] la_oenb[9] la_oenb[8] la_oenb[7] la_oenb[6] la_oenb[5] la_oenb[4]
+ la_oenb[3] la_oenb[2] la_oenb[1] la_oenb[0]
*.iopin vdda1
*.iopin vdda2
*.iopin vssa1
*.iopin vssa2
*.iopin vccd1
*.iopin vccd2
*.iopin vssd1
*.iopin vssd2
*.ipin wb_clk_i
*.ipin wb_rst_i
*.ipin wbs_stb_i
*.ipin wbs_cyc_i
*.ipin wbs_we_i
*.ipin wbs_sel_i[3],wbs_sel_i[2],wbs_sel_i[1],wbs_sel_i[0]
*.ipin
*+ wbs_dat_i[31],wbs_dat_i[30],wbs_dat_i[29],wbs_dat_i[28],wbs_dat_i[27],wbs_dat_i[26],wbs_dat_i[25],wbs_dat_i[24],wbs_dat_i[23],wbs_dat_i[22],wbs_dat_i[21],wbs_dat_i[20],wbs_dat_i[19],wbs_dat_i[18],wbs_dat_i[17],wbs_dat_i[16],wbs_dat_i[15],wbs_dat_i[14],wbs_dat_i[13],wbs_dat_i[12],wbs_dat_i[11],wbs_dat_i[10],wbs_dat_i[9],wbs_dat_i[8],wbs_dat_i[7],wbs_dat_i[6],wbs_dat_i[5],wbs_dat_i[4],wbs_dat_i[3],wbs_dat_i[2],wbs_dat_i[1],wbs_dat_i[0]
*.ipin
*+ wbs_adr_i[31],wbs_adr_i[30],wbs_adr_i[29],wbs_adr_i[28],wbs_adr_i[27],wbs_adr_i[26],wbs_adr_i[25],wbs_adr_i[24],wbs_adr_i[23],wbs_adr_i[22],wbs_adr_i[21],wbs_adr_i[20],wbs_adr_i[19],wbs_adr_i[18],wbs_adr_i[17],wbs_adr_i[16],wbs_adr_i[15],wbs_adr_i[14],wbs_adr_i[13],wbs_adr_i[12],wbs_adr_i[11],wbs_adr_i[10],wbs_adr_i[9],wbs_adr_i[8],wbs_adr_i[7],wbs_adr_i[6],wbs_adr_i[5],wbs_adr_i[4],wbs_adr_i[3],wbs_adr_i[2],wbs_adr_i[1],wbs_adr_i[0]
*.opin wbs_ack_o
*.opin
*+ wbs_dat_o[31],wbs_dat_o[30],wbs_dat_o[29],wbs_dat_o[28],wbs_dat_o[27],wbs_dat_o[26],wbs_dat_o[25],wbs_dat_o[24],wbs_dat_o[23],wbs_dat_o[22],wbs_dat_o[21],wbs_dat_o[20],wbs_dat_o[19],wbs_dat_o[18],wbs_dat_o[17],wbs_dat_o[16],wbs_dat_o[15],wbs_dat_o[14],wbs_dat_o[13],wbs_dat_o[12],wbs_dat_o[11],wbs_dat_o[10],wbs_dat_o[9],wbs_dat_o[8],wbs_dat_o[7],wbs_dat_o[6],wbs_dat_o[5],wbs_dat_o[4],wbs_dat_o[3],wbs_dat_o[2],wbs_dat_o[1],wbs_dat_o[0]
*.ipin
*+ la_data_in[127],la_data_in[126],la_data_in[125],la_data_in[124],la_data_in[123],la_data_in[122],la_data_in[121],la_data_in[120],la_data_in[119],la_data_in[118],la_data_in[117],la_data_in[116],la_data_in[115],la_data_in[114],la_data_in[113],la_data_in[112],la_data_in[111],la_data_in[110],la_data_in[109],la_data_in[108],la_data_in[107],la_data_in[106],la_data_in[105],la_data_in[104],la_data_in[103],la_data_in[102],la_data_in[101],la_data_in[100],la_data_in[99],la_data_in[98],la_data_in[97],la_data_in[96],la_data_in[95],la_data_in[94],la_data_in[93],la_data_in[92],la_data_in[91],la_data_in[90],la_data_in[89],la_data_in[88],la_data_in[87],la_data_in[86],la_data_in[85],la_data_in[84],la_data_in[83],la_data_in[82],la_data_in[81],la_data_in[80],la_data_in[79],la_data_in[78],la_data_in[77],la_data_in[76],la_data_in[75],la_data_in[74],la_data_in[73],la_data_in[72],la_data_in[71],la_data_in[70],la_data_in[69],la_data_in[68],la_data_in[67],la_data_in[66],la_data_in[65],la_data_in[64],la_data_in[63],la_data_in[62],la_data_in[61],la_data_in[60],la_data_in[59],la_data_in[58],la_data_in[57],la_data_in[56],la_data_in[55],la_data_in[54],la_data_in[53],la_data_in[52],la_data_in[51],la_data_in[50],la_data_in[49],la_data_in[48],la_data_in[47],la_data_in[46],la_data_in[45],la_data_in[44],la_data_in[43],la_data_in[42],la_data_in[41],la_data_in[40],la_data_in[39],la_data_in[38],la_data_in[37],la_data_in[36],la_data_in[35],la_data_in[34],la_data_in[33],la_data_in[32],la_data_in[31],la_data_in[30],la_data_in[29],la_data_in[28],la_data_in[27],la_data_in[26],la_data_in[25],la_data_in[24],la_data_in[23],la_data_in[22],la_data_in[21],la_data_in[20],la_data_in[19],la_data_in[18],la_data_in[17],la_data_in[16],la_data_in[15],la_data_in[14],la_data_in[13],la_data_in[12],la_data_in[11],la_data_in[10],la_data_in[9],la_data_in[8],la_data_in[7],la_data_in[6],la_data_in[5],la_data_in[4],la_data_in[3],la_data_in[2],la_data_in[1],la_data_in[0]
*.opin
*+ la_data_out[127],la_data_out[126],la_data_out[125],la_data_out[124],la_data_out[123],la_data_out[122],la_data_out[121],la_data_out[120],la_data_out[119],la_data_out[118],la_data_out[117],la_data_out[116],la_data_out[115],la_data_out[114],la_data_out[113],la_data_out[112],la_data_out[111],la_data_out[110],la_data_out[109],la_data_out[108],la_data_out[107],la_data_out[106],la_data_out[105],la_data_out[104],la_data_out[103],la_data_out[102],la_data_out[101],la_data_out[100],la_data_out[99],la_data_out[98],la_data_out[97],la_data_out[96],la_data_out[95],la_data_out[94],la_data_out[93],la_data_out[92],la_data_out[91],la_data_out[90],la_data_out[89],la_data_out[88],la_data_out[87],la_data_out[86],la_data_out[85],la_data_out[84],la_data_out[83],la_data_out[82],la_data_out[81],la_data_out[80],la_data_out[79],la_data_out[78],la_data_out[77],la_data_out[76],la_data_out[75],la_data_out[74],la_data_out[73],la_data_out[72],la_data_out[71],la_data_out[70],la_data_out[69],la_data_out[68],la_data_out[67],la_data_out[66],la_data_out[65],la_data_out[64],la_data_out[63],la_data_out[62],la_data_out[61],la_data_out[60],la_data_out[59],la_data_out[58],la_data_out[57],la_data_out[56],la_data_out[55],la_data_out[54],la_data_out[53],la_data_out[52],la_data_out[51],la_data_out[50],la_data_out[49],la_data_out[48],la_data_out[47],la_data_out[46],la_data_out[45],la_data_out[44],la_data_out[43],la_data_out[42],la_data_out[41],la_data_out[40],la_data_out[39],la_data_out[38],la_data_out[37],la_data_out[36],la_data_out[35],la_data_out[34],la_data_out[33],la_data_out[32],la_data_out[31],la_data_out[30],la_data_out[29],la_data_out[28],la_data_out[27],la_data_out[26],la_data_out[25],la_data_out[24],la_data_out[23],la_data_out[22],la_data_out[21],la_data_out[20],la_data_out[19],la_data_out[18],la_data_out[17],la_data_out[16],la_data_out[15],la_data_out[14],la_data_out[13],la_data_out[12],la_data_out[11],la_data_out[10],la_data_out[9],la_data_out[8],la_data_out[7],la_data_out[6],la_data_out[5],la_data_out[4],la_data_out[3],la_data_out[2],la_data_out[1],la_data_out[0]
*.ipin
*+ io_in[26],io_in[25],io_in[24],io_in[23],io_in[22],io_in[21],io_in[20],io_in[19],io_in[18],io_in[17],io_in[16],io_in[15],io_in[14],io_in[13],io_in[12],io_in[11],io_in[10],io_in[9],io_in[8],io_in[7],io_in[6],io_in[5],io_in[4],io_in[3],io_in[2],io_in[1],io_in[0]
*.ipin
*+ io_in_3v3[26],io_in_3v3[25],io_in_3v3[24],io_in_3v3[23],io_in_3v3[22],io_in_3v3[21],io_in_3v3[20],io_in_3v3[19],io_in_3v3[18],io_in_3v3[17],io_in_3v3[16],io_in_3v3[15],io_in_3v3[14],io_in_3v3[13],io_in_3v3[12],io_in_3v3[11],io_in_3v3[10],io_in_3v3[9],io_in_3v3[8],io_in_3v3[7],io_in_3v3[6],io_in_3v3[5],io_in_3v3[4],io_in_3v3[3],io_in_3v3[2],io_in_3v3[1],io_in_3v3[0]
*.ipin user_clock2
*.opin
*+ io_out[26],io_out[25],io_out[24],io_out[23],io_out[22],io_out[21],io_out[20],io_out[19],io_out[18],io_out[17],io_out[16],io_out[15],io_out[14],io_out[13],io_out[12],io_out[11],io_out[10],io_out[9],io_out[8],io_out[7],io_out[6],io_out[5],io_out[4],io_out[3],io_out[2],io_out[1],io_out[0]
*.opin
*+ io_oeb[26],io_oeb[25],io_oeb[24],io_oeb[23],io_oeb[22],io_oeb[21],io_oeb[20],io_oeb[19],io_oeb[18],io_oeb[17],io_oeb[16],io_oeb[15],io_oeb[14],io_oeb[13],io_oeb[12],io_oeb[11],io_oeb[10],io_oeb[9],io_oeb[8],io_oeb[7],io_oeb[6],io_oeb[5],io_oeb[4],io_oeb[3],io_oeb[2],io_oeb[1],io_oeb[0]
*.iopin
*+ gpio_analog[17],gpio_analog[16],gpio_analog[15],gpio_analog[14],gpio_analog[13],gpio_analog[12],gpio_analog[11],gpio_analog[10],gpio_analog[9],gpio_analog[8],gpio_analog[7],gpio_analog[6],gpio_analog[5],gpio_analog[4],gpio_analog[3],gpio_analog[2],gpio_analog[1],gpio_analog[0]
*.iopin
*+ gpio_noesd[17],gpio_noesd[16],gpio_noesd[15],gpio_noesd[14],gpio_noesd[13],gpio_noesd[12],gpio_noesd[11],gpio_noesd[10],gpio_noesd[9],gpio_noesd[8],gpio_noesd[7],gpio_noesd[6],gpio_noesd[5],gpio_noesd[4],gpio_noesd[3],gpio_noesd[2],gpio_noesd[1],gpio_noesd[0]
*.iopin
*+ io_analog[10],io_analog[9],io_analog[8],io_analog[7],io_analog[6],io_analog[5],io_analog[4],io_analog[3],io_analog[2],io_analog[1],io_analog[0]
*.iopin io_clamp_high[2],io_clamp_high[1],io_clamp_high[0]
*.iopin io_clamp_low[2],io_clamp_low[1],io_clamp_low[0]
*.opin user_irq[2],user_irq[1],user_irq[0]
*.ipin
*+ la_oenb[127],la_oenb[126],la_oenb[125],la_oenb[124],la_oenb[123],la_oenb[122],la_oenb[121],la_oenb[120],la_oenb[119],la_oenb[118],la_oenb[117],la_oenb[116],la_oenb[115],la_oenb[114],la_oenb[113],la_oenb[112],la_oenb[111],la_oenb[110],la_oenb[109],la_oenb[108],la_oenb[107],la_oenb[106],la_oenb[105],la_oenb[104],la_oenb[103],la_oenb[102],la_oenb[101],la_oenb[100],la_oenb[99],la_oenb[98],la_oenb[97],la_oenb[96],la_oenb[95],la_oenb[94],la_oenb[93],la_oenb[92],la_oenb[91],la_oenb[90],la_oenb[89],la_oenb[88],la_oenb[87],la_oenb[86],la_oenb[85],la_oenb[84],la_oenb[83],la_oenb[82],la_oenb[81],la_oenb[80],la_oenb[79],la_oenb[78],la_oenb[77],la_oenb[76],la_oenb[75],la_oenb[74],la_oenb[73],la_oenb[72],la_oenb[71],la_oenb[70],la_oenb[69],la_oenb[68],la_oenb[67],la_oenb[66],la_oenb[65],la_oenb[64],la_oenb[63],la_oenb[62],la_oenb[61],la_oenb[60],la_oenb[59],la_oenb[58],la_oenb[57],la_oenb[56],la_oenb[55],la_oenb[54],la_oenb[53],la_oenb[52],la_oenb[51],la_oenb[50],la_oenb[49],la_oenb[48],la_oenb[47],la_oenb[46],la_oenb[45],la_oenb[44],la_oenb[43],la_oenb[42],la_oenb[41],la_oenb[40],la_oenb[39],la_oenb[38],la_oenb[37],la_oenb[36],la_oenb[35],la_oenb[34],la_oenb[33],la_oenb[32],la_oenb[31],la_oenb[30],la_oenb[29],la_oenb[28],la_oenb[27],la_oenb[26],la_oenb[25],la_oenb[24],la_oenb[23],la_oenb[22],la_oenb[21],la_oenb[20],la_oenb[19],la_oenb[18],la_oenb[17],la_oenb[16],la_oenb[15],la_oenb[14],la_oenb[13],la_oenb[12],la_oenb[11],la_oenb[10],la_oenb[9],la_oenb[8],la_oenb[7],la_oenb[6],la_oenb[5],la_oenb[4],la_oenb[3],la_oenb[2],la_oenb[1],la_oenb[0]
xtop la_data_in_81_ dvdd gpio_analog_3_ la_data_out_70_ la_data_out_71_ la_data_out_72_
+ la_data_out_73_ la_data_out_74_ la_data_out_75_ la_data_out_76_ la_data_out_77_ la_data_out_78_ la_data_out_79_
+ la_data_out_80_ la_data_in_66_ gpio_analog_2_ la_data_in_82_ avdd la_data_in_69_ vdda1 vssa1 la_data_in_62_ clksys
+ la_data_in_63_ gpio_analog_4_ gpio_analog_5_ la_data_in_67_ la_data_in_68_ la_data_in_61_ gpio_analog_6_
+ la_data_in_42_ la_data_in_43_ la_data_in_44_ avss dvss la_data_in_60_ la_data_in_45_ la_data_in_59_ la_data_in_46_
+ la_data_in_58_ la_data_in_47_ la_data_in_57_ la_data_in_48_ la_data_in_56_ la_data_in_49_ la_data_in_55_
+ la_data_in_50_ la_data_in_54_ la_data_in_51_ la_data_in_53_ la_data_in_52_ top
xsar vdda2 vdda2 vssa2 la_data_out_26_ la_data_out_27_ la_data_out_28_ la_data_out_29_
+ la_data_out_30_ la_data_out_31_ la_data_out_32_ la_data_out_33_ la_data_out_34_ la_data_out_35_ gpio_analog_11_
+ vssa2 gpio_analog_7_ gpio_analog_10_ la_data_in_23_ la_data_out_25_ la_data_in_24_ la_data_in_22_ sar
XC1_447_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_446_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_445_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_444_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_443_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_442_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_441_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_440_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_439_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_438_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_437_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_436_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_435_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_434_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_433_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_432_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_431_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_430_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_429_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_428_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_427_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_426_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_425_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_424_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_423_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_422_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_421_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_420_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_419_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_418_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_417_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_416_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_415_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_414_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_413_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_412_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_411_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_410_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_409_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_408_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_407_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_406_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_405_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_404_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_403_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_402_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_401_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_400_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_399_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_398_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_397_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_396_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_395_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_394_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_393_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_392_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_391_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_390_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_389_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_388_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_387_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_386_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_385_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_384_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_383_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_382_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_381_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_380_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_379_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_378_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_377_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_376_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_375_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_374_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_373_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_372_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_371_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_370_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_369_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_368_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_367_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_366_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_365_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_364_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_363_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_362_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_361_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_360_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_359_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_358_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_357_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_356_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_355_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_354_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_353_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_352_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_351_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_350_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_349_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_348_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_347_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_346_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_345_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_344_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_343_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_342_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_341_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_340_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_339_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_338_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_337_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_336_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_335_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_334_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_333_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_332_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_331_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_330_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_329_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_328_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_327_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_326_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_325_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_324_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_323_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_322_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_321_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_320_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_319_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_318_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_317_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_316_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_315_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_314_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_313_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_312_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_311_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_310_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_309_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_308_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_307_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_306_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_305_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_304_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_303_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_302_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_301_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_300_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_299_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_298_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_297_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_296_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_295_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_294_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_293_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_292_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_291_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_290_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_289_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_288_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_287_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_286_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_285_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_284_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_283_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_282_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_281_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_280_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_279_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_278_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_277_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_276_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_275_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_274_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_273_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_272_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_271_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_270_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_269_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_268_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_267_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_266_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_265_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_264_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_263_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_262_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_261_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_260_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_259_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_258_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_257_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_256_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_255_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_254_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_253_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_252_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_251_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_250_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_249_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_248_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_247_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_246_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_245_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_244_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_243_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_242_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_241_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_240_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_239_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_238_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_237_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_236_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_235_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_234_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_233_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_232_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_231_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_230_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_229_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_228_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_227_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_226_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_225_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_224_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_223_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_222_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_221_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_220_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_219_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_218_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_217_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_216_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_215_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_214_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_213_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_212_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_211_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_210_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_209_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_208_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_207_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_206_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_205_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_204_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_203_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_202_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_201_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_200_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_199_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_198_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_197_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_196_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_195_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_194_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_193_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_192_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_191_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_190_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_189_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_188_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_187_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_186_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_185_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_184_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_183_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_182_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_181_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_180_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_179_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_178_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_177_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_176_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_175_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_174_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_173_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_172_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_171_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_170_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_169_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_168_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_167_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_166_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_165_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_164_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_163_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_162_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_161_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_160_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_159_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_158_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_157_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_156_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_155_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_154_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_153_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_152_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_151_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_150_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_149_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_148_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_147_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_146_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_145_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_144_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_143_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_142_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_141_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_140_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_139_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_138_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_137_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_136_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_135_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_134_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_133_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_132_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_131_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_130_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_129_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_128_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_127_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_126_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_125_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_124_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_123_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_122_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_121_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_120_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_119_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_118_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_117_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_116_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_115_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_114_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_113_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_112_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_111_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_110_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_109_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_108_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_107_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_106_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_105_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_104_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_103_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_102_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_101_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_100_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_99_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_98_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_97_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_96_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_95_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_94_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_93_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_92_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_91_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_90_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_89_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_88_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_87_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_86_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_85_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_84_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_83_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_82_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_81_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_80_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_79_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_78_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_77_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_76_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_75_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_74_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_73_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_72_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_71_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_70_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_69_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_68_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_67_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_66_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_65_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_64_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_63_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_62_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_61_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_60_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_59_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_58_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_57_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_56_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_55_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_54_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_53_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_52_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_51_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_50_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_49_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_48_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_47_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_46_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_45_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_44_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_43_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_42_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_41_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_40_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_39_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_38_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_37_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_36_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_35_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_34_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_33_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_32_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_31_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_30_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_29_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_28_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_27_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_26_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_25_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_24_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_23_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_22_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_21_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_20_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_19_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_18_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_17_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_16_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_15_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_14_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_13_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_12_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_11_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_10_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_9_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_8_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_7_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_6_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_5_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_4_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_3_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_2_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_1_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
XC1_0_ vdda2 vssa2 sky130_fd_pr__cap_mim_m3_2 W=30 L=30 MF=1 m=1
.ends


* expanding   symbol:  top/top.sym # of pins=25
* sym_path: /home/christoph/Studium/projekte/design/design/top/top.sym
* sch_path: /home/christoph/Studium/projekte/design/design/top/top.sch
.subckt top  en_caladc dvdd inp result_9_ result_8_ result_7_ result_6_ result_5_ result_4_
+ result_3_ result_2_ result_1_ result_0_ valid en_ldo_dig inn en_adc avdd rstn vdd vss en_ldo_ana clksys
+ en_clk_int clkext tbout en_clkdiv clksel refsel vbg_ext tbctl_2_ tbctl_1_ tbctl_0_ avss dvss bgtrim_15_
+ bgtrim_14_ bgtrim_13_ bgtrim_12_ bgtrim_11_ bgtrim_10_ bgtrim_9_ bgtrim_8_ bgtrim_7_ bgtrim_6_ bgtrim_5_
+ bgtrim_4_ bgtrim_3_ bgtrim_2_ bgtrim_1_ bgtrim_0_
*.ipin inp
*.ipin inn
*.ipin clksel
*.ipin clkext
*.ipin en_caladc
*.ipin en_adc
*.ipin en_clkdiv
*.opin clksys
*.ipin en_ldo_ana
*.ipin en_ldo_dig
*.opin
*+ result_9_,result_8_,result_7_,result_6_,result_5_,result_4_,result_3_,result_2_,result_1_,result_0_
*.opin valid
*.ipin refsel
*.iopin vdd
*.iopin vss
*.ipin rstn
*.ipin vbg_ext
*.ipin en_clk_int
*.iopin avdd
*.iopin dvdd
*.opin tbout
*.iopin avss
*.iopin dvss
*.ipin
*+ bgtrim_15_,bgtrim_14_,bgtrim_13_,bgtrim_12_,bgtrim_11_,bgtrim_10_,bgtrim_9_,bgtrim_8_,bgtrim_7_,bgtrim_6_,bgtrim_5_,bgtrim_4_,bgtrim_3_,bgtrim_2_,bgtrim_1_,bgtrim_0_
*.ipin tbctl_2_,tbctl_1_,tbctl_0_
xm dvdd en_ldo_dig avdd rstn vdd vss en_ldo_ana clksys en_clk_int clkext ibp_3_ ibp_2_ ibp_1_ ibp_0_
+ ibn_1_ ibn_0_ en_clkdiv clksel refsel vbg_ext avss dvss tbout bgtrim_15_ bgtrim_14_ bgtrim_13_ bgtrim_12_
+ bgtrim_11_ bgtrim_10_ bgtrim_9_ bgtrim_8_ bgtrim_7_ bgtrim_6_ bgtrim_5_ bgtrim_4_ bgtrim_3_ bgtrim_2_
+ bgtrim_1_ bgtrim_0_ tbctl_2_ tbctl_1_ tbctl_0_ main
xsar avdd dvdd dvss result_9_ result_8_ result_7_ result_6_ result_5_ result_4_ result_3_ result_2_
+ result_1_ result_0_ inn avss clksys inp en_adc valid en_caladc rstn sar
.ends


* expanding   symbol:  sar_10b/sar/sar.sym # of pins=12
* sym_path: /home/christoph/Studium/projekte/design/design/sar_10b/sar/sar.sym
* sch_path: /home/christoph/Studium/projekte/design/design/sar_10b/sar/sar.sch
.subckt sar  avdd dvdd dvss result_9_ result_8_ result_7_ result_6_ result_5_ result_4_ result_3_
+ result_2_ result_1_ result_0_ vinn avss clk vinp en valid cal rstn
*.iopin avss
*.iopin avdd
*.iopin dvss
*.iopin dvdd
*.ipin vinp
*.ipin vinn
*.opin
*+ result_9_,result_8_,result_7_,result_6_,result_5_,result_4_,result_3_,result_2_,result_1_,result_0_
*.ipin clk
*.ipin en
*.opin valid
*.ipin cal
*.ipin rstn
xlat dvdd comp net1 dvss outn outp latch
xdn vn sample avdd avss vinn ctln_9_ ctln_8_ ctln_7_ ctln_6_ ctln_5_ ctln_4_ ctln_3_ ctln_2_ ctln_1_
+ ctln_0_ avss dac
xdp vp sample avdd avss vinp ctlp_9_ ctlp_8_ ctlp_7_ ctlp_6_ ctlp_5_ ctlp_4_ ctlp_3_ ctlp_2_ ctlp_1_
+ ctlp_0_ avdd dac
xcom avss avdd clkca outp vp outn vn trim_4_ trim_3_ trim_2_ trim_1_ trim_0_ trimb_4_ trimb_3_
+ trimb_2_ trimb_1_ trimb_0_ comparator
XC1_57_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_56_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_55_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_54_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_53_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_52_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_51_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_50_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_49_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_48_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_47_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_46_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_45_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_44_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_43_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_42_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_41_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_40_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_39_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_38_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_37_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_36_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_35_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_34_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_33_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_32_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_31_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_30_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_29_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_28_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_27_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_26_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_25_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_24_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_23_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_22_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_21_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_20_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_19_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_18_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_17_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_16_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_15_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_14_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_13_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_12_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_11_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_10_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_9_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_8_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_7_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_6_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_5_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_4_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_3_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_2_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_1_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC1_0_ avdd avss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC2_13_ dvdd dvss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC2_12_ dvdd dvss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC2_11_ dvdd dvss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC2_10_ dvdd dvss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC2_9_ dvdd dvss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC2_8_ dvdd dvss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC2_7_ dvdd dvss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC2_6_ dvdd dvss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC2_5_ dvdd dvss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC2_4_ dvdd dvss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC2_3_ dvdd dvss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC2_2_ dvdd dvss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC2_1_ dvdd dvss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
XC2_0_ dvdd dvss sky130_fd_pr__cap_mim_m3_2 W=12 L=12 MF=1 m=1
xlogic trim_4_ trim_3_ trim_2_ trim_1_ trim_0_ trimb_4_ trimb_3_ trimb_2_ trimb_1_ trimb_0_ clkc
+ comp cal en ctlp_9_ ctlp_8_ ctlp_7_ ctlp_6_ ctlp_5_ ctlp_4_ ctlp_3_ ctlp_2_ ctlp_1_ ctlp_0_ clk
+ result_9_ result_8_ result_7_ result_6_ result_5_ result_4_ result_3_ result_2_ result_1_ result_0_ ctln_9_
+ ctln_8_ ctln_7_ ctln_6_ ctln_5_ ctln_4_ ctln_3_ ctln_2_ ctln_1_ ctln_0_ valid rstn sample dvdd dvss
+ sarlogic
xbuf avdd clkc clkca avss buffer_lvt
.ends


* expanding   symbol:  main/main.sym # of pins=21
* sym_path: /home/christoph/Studium/projekte/design/design/main/main.sym
* sch_path: /home/christoph/Studium/projekte/design/design/main/main.sch
.subckt main  dvdd en_ldo_dig avdd rstn vdd vss en_ldo_ana clksys en_clk_int clkext ibp_3_ ibp_2_
+ ibp_1_ ibp_0_ ibn_1_ ibn_0_ en_clkdiv clksel refsel vbg_ext avss dvss tbout bgtrim_15_ bgtrim_14_
+ bgtrim_13_ bgtrim_12_ bgtrim_11_ bgtrim_10_ bgtrim_9_ bgtrim_8_ bgtrim_7_ bgtrim_6_ bgtrim_5_ bgtrim_4_
+ bgtrim_3_ bgtrim_2_ bgtrim_1_ bgtrim_0_ tbctl_2_ tbctl_1_ tbctl_0_
*.ipin clksel
*.ipin clkext
*.ipin en_clkdiv
*.ipin en_ldo_ana
*.ipin en_ldo_dig
*.ipin en_clk_int
*.ipin vbg_ext
*.ipin refsel
*.opin ibp_3_,ibp_2_,ibp_1_,ibp_0_
*.opin ibn_1_,ibn_0_
*.iopin vdd
*.iopin vss
*.ipin rstn
*.opin clksys
*.iopin dvss
*.iopin avss
*.iopin dvdd
*.iopin avdd
*.ipin
*+ bgtrim_15_,bgtrim_14_,bgtrim_13_,bgtrim_12_,bgtrim_11_,bgtrim_10_,bgtrim_9_,bgtrim_8_,bgtrim_7_,bgtrim_6_,bgtrim_5_,bgtrim_4_,bgtrim_3_,bgtrim_2_,bgtrim_1_,bgtrim_0_
*.opin tbout
*.ipin tbctl_2_,tbctl_1_,tbctl_0_
xbg vdd vbg_int vss ibnbas bgtrim_15_ bgtrim_14_ bgtrim_13_ bgtrim_12_ bgtrim_11_ bgtrim_10_
+ bgtrim_9_ bgtrim_8_ bgtrim_7_ bgtrim_6_ bgtrim_5_ bgtrim_4_ bgtrim_3_ bgtrim_2_ bgtrim_1_ bgtrim_0_ bandgap
xbb ibpbas vbg ibp_3_ ibp_2_ ibp_1_ ibp_0_ ibn_1_ ibn_0_ vdd vss vb_6_ vb_5_ vb_4_ vb_3_ vb_2_ vb_1_
+ vb_0_ bias
xro avdd avss dvdd dvss rstn ibn_0_ clkint en_clk_int rosc
xbc vdd vss ibpbas ibnbas bias_basis_current
xra avdd vb_2_ vss vdd ibp_1_ en_ldo_ana avdd regulator
xrd dvdd vb_3_ vss vdd ibp_2_ en_ldo_dig dvdd regulator
xcs dvdd dvss rstn clkint clksys clkext en_clkdiv clksel clksel
xsw vbg refsel vdd vbg_ext vss vbg_int spdt
xtb ibp_0_ tbout vdd vss vbg vss dvdd vb_4_ vb_3_ vb_2_ avdd tbctl_2_ tbctl_1_ tbctl_0_ testbuffer
R3 vss avss sky130_fd_pr__res_generic_m4 W=9.6 L=4 m=1
R1 vss dvss sky130_fd_pr__res_generic_m4 W=9.6 L=4 m=1
.ends


* expanding   symbol:  sar_10b/latch/latch.sym # of pins=6
* sym_path: /home/christoph/Studium/projekte/design/design/sar_10b/latch/latch.sym
* sch_path: /home/christoph/Studium/projekte/design/design/sar_10b/latch/latch.sch
.subckt latch  vdd Q Qn vss R S
*.ipin S
*.ipin R
*.iopin vss
*.iopin vdd
*.opin Q
*.opin Qn
x1 vdd Qn Q vss inv_lvt
x2 vdd Q Qn vss inv_lvt
x3 vdd R net2 vss inv_lvt
x4 vdd S net1 vss inv_lvt
XM3 Qn net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 Q net2 vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  sar_10b/dac/dac.sym # of pins=7
* sym_path: /home/christoph/Studium/projekte/design/design/sar_10b/dac/dac.sym
* sch_path: /home/christoph/Studium/projekte/design/design/sar_10b/dac/dac.sch
.subckt dac  out sample vdd vss vin ctl_9_ ctl_8_ ctl_7_ ctl_6_ ctl_5_ ctl_4_ ctl_3_ ctl_2_ ctl_1_
+ ctl_0_ dum
*.ipin vin
*.ipin sample
*.opin out
*.ipin ctl_9_,ctl_8_,ctl_7_,ctl_6_,ctl_5_,ctl_4_,ctl_3_,ctl_2_,ctl_1_,ctl_0_
*.ipin dum
*.iopin vdd
*.iopin vss
xca out n6 n0 n5 n4 n2 ndum n3 n1 n7 n8 n9 carray
xswt out sample vdd vin vss bootstrapped_sw_hv
xidum dum vss vss vdd vdd ndum sky130_fd_sc_hd__inv_2
xi0 ctl_0_ vss vss vdd vdd n0 sky130_fd_sc_hd__inv_2
xi1 ctl_1_ vss vss vdd vdd n1 sky130_fd_sc_hd__inv_2
xi2 ctl_2_ vss vss vdd vdd n2 sky130_fd_sc_hd__inv_2
xi3 ctl_3_ vss vss vdd vdd n3 sky130_fd_sc_hd__inv_2
xi4 ctl_4_ vss vss vdd vdd n4 sky130_fd_sc_hd__inv_2
xi5 ctl_5_ vss vss vdd vdd n5 sky130_fd_sc_hd__inv_2
xi6 ctl_6_ vss vss vdd vdd n6 sky130_fd_sc_hd__inv_2
xi7 ctl_7_ vss vss vdd vdd n7 sky130_fd_sc_hd__inv_2
xi8 ctl_8_ vss vss vdd vdd n8 sky130_fd_sc_hd__inv_2
xi9 ctl_9_ vss vss vdd vdd n9 sky130_fd_sc_hd__inv_2
.ends


* expanding   symbol:  sar_10b/comparator/comparator.sym # of pins=9
* sym_path: /home/christoph/Studium/projekte/design/design/sar_10b/comparator/comparator.sym
* sch_path: /home/christoph/Studium/projekte/design/design/sar_10b/comparator/comparator.sch
.subckt comparator  vss vdd clk outp vp outn vn trim_4_ trim_3_ trim_2_ trim_1_ trim_0_ trimb_4_
+ trimb_3_ trimb_2_ trimb_1_ trimb_0_
*.ipin vn
*.ipin vp
*.ipin clk
*.iopin vdd
*.iopin vss
*.opin outp
*.opin outn
*.ipin trim_4_,trim_3_,trim_2_,trim_1_,trim_0_
*.ipin trimb_4_,trimb_3_,trimb_2_,trimb_1_,trimb_0_
XMdiff diff clk vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XMinn in vn diff vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMinp ip vp diff vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMl4 outp outn vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMl3 outn outp vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 outp clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 outn clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMl1 outn outp in vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMl2 outp outn ip vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 ip clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 in clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
x2 in trim_4_ trim_3_ trim_2_ trim_1_ trim_0_ vss trim
x3 ip trimb_4_ trimb_3_ trimb_2_ trimb_1_ trimb_0_ vss trim
.ends


* expanding   symbol:  sar_10b/control/sarlogic.sym # of pins=15
* sym_path: /home/christoph/Studium/projekte/design/design/sar_10b/control/sarlogic.sym
* sch_path: /home/christoph/Studium/projekte/design/design/sar_10b/control/sarlogic.sch
.subckt sarlogic  trim_4_ trim_3_ trim_2_ trim_1_ trim_0_ trimb_4_ trimb_3_ trimb_2_ trimb_1_
+ trimb_0_ clkc comp cal en ctlp_9_ ctlp_8_ ctlp_7_ ctlp_6_ ctlp_5_ ctlp_4_ ctlp_3_ ctlp_2_ ctlp_1_ ctlp_0_
+ clk result_9_ result_8_ result_7_ result_6_ result_5_ result_4_ result_3_ result_2_ result_1_ result_0_
+ ctln_9_ ctln_8_ ctln_7_ ctln_6_ ctln_5_ ctln_4_ ctln_3_ ctln_2_ ctln_1_ ctln_0_ valid rstn sample dvdd dvss
*.opin clkc
*.opin ctlp_9_,ctlp_8_,ctlp_7_,ctlp_6_,ctlp_5_,ctlp_4_,ctlp_3_,ctlp_2_,ctlp_1_,ctlp_0_
*.opin ctln_9_,ctln_8_,ctln_7_,ctln_6_,ctln_5_,ctln_4_,ctln_3_,ctln_2_,ctln_1_,ctln_0_
*.opin sample
*.opin trim_4_,trim_3_,trim_2_,trim_1_,trim_0_
*.opin trimb_4_,trimb_3_,trimb_2_,trimb_1_,trimb_0_
*.ipin comp
*.ipin cal
*.ipin en
*.ipin clk
*.ipin
*+ result_9_,result_8_,result_7_,result_6_,result_5_,result_4_,result_3_,result_2_,result_1_,result_0_
*.ipin rstn
*.iopin dvdd
*.iopin dvss
*.opin valid
**** begin user architecture code
.include /home/christoph/Studium/projekte/design/design/sar_10b/control/cmos_cells_digital.sp
.include /home/christoph/Studium/projekte/design/design/sar_10b/control/sarlogic.sp

**** end user architecture code
**** begin user architecture code
* Keep the sar_logic underscore name. Otherwise xschem gets confused.
Xuut dclk drstn den dcomp dcal dvalid dres0 dres1 dres2 dres3 dres4 dres5 dres6 dres7 dres8 dres9
+ dsamp dctlp0 dctlp1 dctlp2 dctlp3 dctlp4 dctlp5 dctlp6 dctlp7 dctlp8 dctlp9 dctln0 dctln1 dctln2 dctln3
+ dctln4 dctln5 dctln6 dctln7 dctln8 dctln9 dtrim0 dtrim1 dtrim2 dtrim3 dtrim4 dtrimb0 dtrimb1 dtrimb2
+ dtrimb3 dtrimb4 dclkc sar_logic

.model adc_buff adc_bridge(in_low = 0.2 in_high=0.8)
.model dac_buff dac_bridge(out_high = 1.2)

Aad [clk rstn en comp cal] [dclk drstn den dcomp dcal] adc_buff
Ada1 [dctlp0 dctlp1 dctlp2 dctlp3 dctlp4 dctlp5 dctlp6 dctlp7 dctlp8 dctlp9] [ctlp_0_ ctlp_1_
+ ctlp_2_ ctlp_3_ ctlp_4_ ctlp_5_ ctlp_6_ ctlp_7_ ctlp_8_ ctlp_9_] dac_buff
Ada2 [dctln0 dctln1 dctln2 dctln3 dctln4 dctln5 dctln6 dctln7 dctln8 dctln9] [ctln_0_ ctln_1_
+ ctln_2_ ctln_3_ ctln_4_ ctln_5_ ctln_6_ ctln_7_ ctln_8_ ctln_9_] dac_buff
Ada3 [dres0 dres1 dres2 dres3 dres4 dres5 dres6 dres7 dres8 dres9 dsamp dclkc] [res0 res1 res2 res3
+ res4 res5 res6 res7 res8 res9 sample clkc] dac_buff
Ada4 [dtrim4 dtrim3 dtrim2 dtrim1 dtrim0 dtrimb4 dtrimb3 dtrimb2 dtrimb1 dtrimb0] [trim_4_ trim_3_
+ trim_2_ trim_1_ trim_0_ trimb_4_ trimb_3_ trimb_2_ trimb_1_ trimb_0_ ] dac_buff
Ada5 [dvalid] [valid] dac_buff

**** end user architecture code
.ends


* expanding   symbol:  logic/buffer_lvt.sym # of pins=4
* sym_path: /home/christoph/Studium/projekte/design/design/logic/buffer_lvt.sym
* sch_path: /home/christoph/Studium/projekte/design/design/logic/buffer_lvt.sch
.subckt buffer_lvt  vdd in out vss
*.iopin vdd
*.iopin vss
*.ipin in
*.opin out
XM1 net1 in vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 net1 in vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 out net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 out net1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  bandgap/bandgap.sym # of pins=5
* sym_path: /home/christoph/Studium/projekte/design/design/bandgap/bandgap.sym
* sch_path: /home/christoph/Studium/projekte/design/design/bandgap/bandgap.sch
.subckt bandgap  vdd vbg vss bias trim_15_ trim_14_ trim_13_ trim_12_ trim_11_ trim_10_ trim_9_
+ trim_8_ trim_7_ trim_6_ trim_5_ trim_4_ trim_3_ trim_2_ trim_1_ trim_0_
*.iopin vdd
*.iopin vss
*.opin vbg
*.iopin bias
*.ipin
*+ trim_15_,trim_14_,trim_13_,trim_12_,trim_11_,trim_10_,trim_9_,trim_8_,trim_7_,trim_6_,trim_5_,trim_4_,trim_3_,trim_2_,trim_1_,trim_0_
XQ2 vss vss em2 vss sky130_fd_pr__pnp_05v5_W0p68L0p68 m=8
XQ1 vss vss vn vss sky130_fd_pr__pnp_05v5_W0p68L0p68 m=1
XC1 gate vss sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=8 m=8
xres vbg comp vp vn vss bg_res
XR1 net1 vp vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XM1 comp gate vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM2 vbg gate vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
xtr net1 em2 trim_15_ trim_14_ trim_13_ trim_12_ trim_11_ trim_10_ trim_9_ trim_8_ trim_7_ trim_6_
+ trim_5_ trim_4_ trim_3_ trim_2_ trim_1_ trim_0_ vss bg_trim
xamp vdd gate vp vn vss bias se_folded_cascode_p
XM3 vs1 vbg vss vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 gate vs1 vss vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 vs1 vs2 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XC2 vs2 vss sky130_fd_pr__cap_mim_m3_1 W=10 L=10 MF=3 m=3
XM6 vs2 vs2 vdd vdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7 vss vdd vs2 vs2 sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  bias/bias.sym # of pins=7
* sym_path: /home/christoph/Studium/projekte/design/design/bias/bias.sym
* sch_path: /home/christoph/Studium/projekte/design/design/bias/bias.sch
.subckt bias  iamp vbg ibp_3_ ibp_2_ ibp_1_ ibp_0_ ibn_1_ ibn_0_ vdd vss vb_6_ vb_5_ vb_4_ vb_3_
+ vb_2_ vb_1_ vb_0_
*.ipin vbg
*.ipin iamp
*.iopin vdd
*.iopin ibp_3_,ibp_2_,ibp_1_,ibp_0_
*.iopin ibn_1_,ibn_0_
*.iopin vb_6_,vb_5_,vb_4_,vb_3_,vb_2_,vb_1_,vb_0_
*.iopin vss
x1 vdd gate fb vbg vss iamp bias_amp
XMP2_1_ gate_cas gate net1_1_ vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMP2_0_ gate_cas gate net1_0_ vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM1 fb gate vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XMPS2_1_ net1_1_ gate vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMPS2_0_ net1_0_ gate vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMP4_1_ ibp_1_ gate net2_1_ vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMP4_0_ ibp_1_ gate net2_0_ vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMPS4_1_ net2_1_ gate vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMPS4_0_ net2_0_ gate vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMP5_1_ ibp_2_ gate net3_1_ vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMP5_0_ ibp_2_ gate net3_0_ vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMPS5_1_ net3_1_ gate vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMPS5_0_ net3_0_ gate vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMP6_1_ ibp_3_ gate net4_1_ vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMP6_0_ ibp_3_ gate net4_0_ vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMPS6_1_ net4_1_ gate vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMPS6_0_ net4_0_ gate vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMP3_3_ ibp_0_ gate net5_3_ vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMP3_2_ ibp_0_ gate net5_2_ vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMP3_1_ ibp_0_ gate net5_1_ vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMP3_0_ ibp_0_ gate net5_0_ vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMPS3_3_ net5_3_ gate vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMPS3_2_ net5_2_ gate vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMPS3_1_ net5_1_ gate vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMPS3_0_ net5_0_ gate vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMNS2_3_ gate_n gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMNS2_2_ gate_n gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMNS2_1_ gate_n gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMNS2_0_ gate_n gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMNS3_3_ net6_3_ gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMNS3_2_ net6_2_ gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMNS3_1_ net6_1_ gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMNS3_0_ net6_0_ gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMNS4_3_ net7_3_ gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMNS4_2_ net7_2_ gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMNS4_1_ net7_1_ gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMNS4_0_ net7_0_ gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMN2_3_ gate_cas gate_cas gate_n vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMN2_2_ gate_cas gate_cas gate_n vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMN2_1_ gate_cas gate_cas gate_n vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMN2_0_ gate_cas gate_cas gate_n vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMN3_3_ ibn_0_ gate_cas net6_3_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMN3_2_ ibn_0_ gate_cas net6_2_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMN3_1_ ibn_0_ gate_cas net6_1_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMN3_0_ ibn_0_ gate_cas net6_0_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMN4_3_ ibn_1_ gate_cas net7_3_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMN4_2_ ibn_1_ gate_cas net7_2_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMN4_1_ ibn_1_ gate_cas net7_1_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMN4_0_ ibn_1_ gate_cas net7_0_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XC1 gate fb sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=8 m=8
XR1 fb net8 vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR2 net8 vb_0_ vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR3 vb_0_ net9 vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR4 net9 vb_1_ vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR5 vb_2_ net11 vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR6 net11 vb_1_ vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR7 vb_3_ net10 vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR8 net10 vb_2_ vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR9 vb_3_ net12 vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR10 net12 vb_4_ vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR11 vb_4_ net13 vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR12 net13 vb_5_ vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR13 vb_6_ net15 vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR14 net15 vb_5_ vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR15 vss net14 vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR16 net14 vb_6_ vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XMP1 vdd gate vdd vdd sky130_fd_pr__pfet_01v8_lvt L=2 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=24 m=24 
XMDUM_7_ vss gate_cas vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM_6_ vss gate_cas vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM_5_ vss gate_cas vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM_4_ vss gate_cas vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM_3_ vss gate_cas vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM_2_ vss gate_cas vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM_1_ vss gate_cas vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM_0_ vss gate_cas vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM_1_3_ vss gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM_1_2_ vss gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM_1_1_ vss gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM_1_0_ vss gate_n vss vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_3_ ibn_0_ gate_cas ibn_0_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_2_ ibn_0_ gate_cas ibn_0_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_1_ ibn_0_ gate_cas ibn_0_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_0_ ibn_0_ gate_cas ibn_0_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_3_ ibn_1_ gate_cas ibn_1_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_2_ ibn_1_ gate_cas ibn_1_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_1_ ibn_1_ gate_cas ibn_1_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_0_ ibn_1_ gate_cas ibn_1_ vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_3_ gate_cas gate_cas gate_cas vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_2_ gate_cas gate_cas gate_cas vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_1_ gate_cas gate_cas gate_cas vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_0_ gate_cas gate_cas gate_cas vss sky130_fd_pr__nfet_01v8_lvt L=2 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XR17_1_ vss vss vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
XR17_0_ vss vss vss sky130_fd_pr__res_xhigh_po W=0.69 L=25.8 mult=1 m=1
.ends


* expanding   symbol:  rosc/rosc.sym # of pins=8
* sym_path: /home/christoph/Studium/projekte/design/design/rosc/rosc.sym
* sch_path: /home/christoph/Studium/projekte/design/design/rosc/rosc.sch
.subckt rosc  avdd avss dvdd dvss rst_b ibias clk en
*.ipin en
*.iopin avss
*.opin clk
*.iopin dvdd
*.iopin dvss
*.iopin avdd
*.ipin rst_b
*.ipin ibias
x8 clk dvss dvss dvdd dvdd fb sky130_fd_sc_hd__inv_1
XM2 bias_n ibias avdd avdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM1 ibias ibias avdd avdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
x9 out_dig fb rst_b dvss dvss dvdd dvdd clk net2 sky130_fd_sc_hd__dfrbp_2
XM4 bias_n bias_n avss avss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM5 vn bias_n avss avss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
x7 out_ana dvss dvss dvdd dvdd out_dig sky130_fd_sc_hd__inv_1
XM3 vp ibias avdd avdd sky130_fd_pr__pfet_01v8 L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XC1 out1 avss sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1 m=1
XC2 out2 avss sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1 m=1
x6 avdd out7 out_ana avss inv_lvt
XM6 out2 out1 vn avss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7 out2 out1 vp avdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XC3 out3 avss sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1 m=1
XC4 out4 avss sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1 m=1
XC5 out5 avss sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1 m=1
XC6 out6 avss sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1 m=1
XM18 net1 out7 vn avss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM19 out1 en vp avdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM20 out1 en net1 avss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM21 out1 out7 vp avdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM8 out3 out2 vn avss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM9 out3 out2 vp avdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM10 out4 out3 vn avss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM11 out4 out3 vp avdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM12 out5 out4 vn avss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM13 out5 out4 vp avdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM14 out6 out5 vn avss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM15 out6 out5 vp avdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM16 out7 out6 vn avss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM17 out7 out6 vp avdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XC7 out7 avss sky130_fd_pr__cap_mim_m3_1 W=4 L=4 MF=1 m=1
.ends


* expanding   symbol:  bias/bias_basis_current.sym # of pins=4
* sym_path: /home/christoph/Studium/projekte/design/design/bias/bias_basis_current.sym
* sch_path: /home/christoph/Studium/projekte/design/design/bias/bias_basis_current.sch
.subckt bias_basis_current  vdd vss ibp ibn
*.iopin ibn
*.iopin vdd
*.iopin vss
*.iopin ibp
XM5 vbp vbp vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM4 vbn vbp vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM1 vbn vbn vss vss sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM2 vbp vbn vres vss sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=32 m=32 
XM6 ibp vbp vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM3 ibn vbn vss vss sky130_fd_pr__nfet_01v8_lvt L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM7 vsu vsu vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM8 vdd vsu vbn vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM9 vsu vsu net1 vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM10 net1 net1 net2 vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XR2 vss vres vss sky130_fd_pr__res_xhigh_po W=0.35 L=14 mult=1 m=1
XR1 net2 vdd vss sky130_fd_pr__res_xhigh_po W=0.35 L=17 mult=1 m=1
.ends


* expanding   symbol:  regulator/regulator.sym # of pins=7
* sym_path: /home/christoph/Studium/projekte/design/design/regulator/regulator.sym
* sch_path: /home/christoph/Studium/projekte/design/design/regulator/regulator.sch
.subckt regulator  out vref vss vin bias en fb
*.iopin vin
*.iopin vss
*.ipin vref
*.opin out
*.iopin bias
*.ipin en
*.ipin fb
XM2 comp vref diff vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM1 mirr fbdiv diff vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM5 diff bias vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM4 comp mirr vin vin sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM3 mirr mirr vin vin sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM6 bias bias vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM7_31_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_30_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_29_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_28_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_27_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_26_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_25_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_24_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_23_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_22_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_21_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_20_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_19_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_18_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_17_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_16_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_15_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_14_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_13_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_12_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_11_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_10_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XM7_9_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7_8_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7_7_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7_6_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7_5_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7_4_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7_3_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7_2_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7_1_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7_0_ out comp vin vin sky130_fd_pr__pfet_01v8_lvt L=0.5 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XC1 out comp sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=8 m=8
XM9 bias enb vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
x1 vin en enb vss inv_lvt
XM8 comp en vin vin sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM10 bias bias bias vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM11 diff bias diff vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM12 comp comp comp vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM13 mirr mirr mirr vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM15 mirr mirr mirr vin sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XM16 comp mirr comp vin sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=2 m=2 
XR2 fbdiv fb vss sky130_fd_pr__res_xhigh_po W=0.35 L=34 mult=1 m=1
XR1 vss fbdiv vss sky130_fd_pr__res_xhigh_po W=0.35 L=34 mult=1 m=1
XR3_1_ vss vss vss sky130_fd_pr__res_xhigh_po W=0.35 L=8.5 mult=1 m=1
XR3_0_ vss vss vss sky130_fd_pr__res_xhigh_po W=0.35 L=8.5 mult=1 m=1
.ends


* expanding   symbol:  clksel/clksel.sym # of pins=8
* sym_path: /home/christoph/Studium/projekte/design/design/clksel/clksel.sym
* sch_path: /home/christoph/Studium/projekte/design/design/clksel/clksel.sch
.subckt clksel  dvdd dvss rst_b clk_int clk_out clk_ext en_div clk_sel
*.ipin clk_int
*.ipin rst_b
*.opin clk_out
*.iopin dvdd
*.iopin dvss
*.ipin clk_ext
*.ipin en_div
*.ipin clk_sel
x1 dvss net2 net3 rst_b dvdd clkdiv
x2 clk_int clk_ext clk_sel dvss dvss dvdd dvdd net2 sky130_fd_sc_hd__mux2_2
x3 net1 dvss dvss dvdd dvdd clk_out sky130_fd_sc_hd__clkbuf_8
x4 net2 net3 en_div dvss dvss dvdd dvdd net1 sky130_fd_sc_hd__mux2_2
.ends


* expanding   symbol:  support/spdt.sym # of pins=6
* sym_path: /home/christoph/Studium/projekte/design/design/support/spdt.sym
* sch_path: /home/christoph/Studium/projekte/design/design/support/spdt.sch
.subckt spdt  out en vdd inb vss ina
*.ipin en
*.iopin vss
*.iopin vdd
*.iopin ina
*.iopin out
*.iopin inb
xinv vdd en enb vss inv_lvt
xsa out en vdd ina vss passgate
xsb out enb vdd inb vss passgate
.ends


* expanding   symbol:  testbuffer/testbuffer.sym # of pins=6
* sym_path: /home/christoph/Studium/projekte/design/design/testbuffer/testbuffer.sym
* sch_path: /home/christoph/Studium/projekte/design/design/testbuffer/testbuffer.sch
.subckt testbuffer  bias out vdd vss inp_6_ inp_5_ inp_4_ inp_3_ inp_2_ inp_1_ inp_0_ ctl_2_ ctl_1_
+ ctl_0_
*.iopin out
*.iopin vss
*.iopin vdd
*.iopin bias
*.ipin inp_6_,inp_5_,inp_4_,inp_3_,inp_2_,inp_1_,inp_0_
*.ipin ctl_2_,ctl_1_,ctl_0_
xmux mux_out vdd vss inp_6_ inp_5_ inp_4_ inp_3_ inp_2_ inp_1_ inp_0_ vdd ctl_2_ ctl_1_ ctl_0_ mux
xamp vdd out mux_out out vss bias se_folded_cascode_np_ab
.ends


* expanding   symbol:  logic/inv_lvt.sym # of pins=4
* sym_path: /home/christoph/Studium/projekte/design/design/logic/inv_lvt.sym
* sch_path: /home/christoph/Studium/projekte/design/design/logic/inv_lvt.sch
.subckt inv_lvt  vdd in out vss
*.iopin vdd
*.iopin vss
*.ipin in
*.opin out
XM1 out in vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  sar_10b/dac/carray.sym # of pins=12
* sym_path: /home/christoph/Studium/projekte/design/design/sar_10b/dac/carray.sym
* sch_path: /home/christoph/Studium/projekte/design/design/sar_10b/dac/carray.sch
.subckt carray  top n6 n0 n5 n4 n2 ndum n3 n1 n7 n8 n9
*.iopin top
*.iopin n7
*.iopin n6
*.iopin n5
*.iopin n4
*.iopin n2
*.iopin n0
*.iopin ndum
*.iopin n3
*.iopin n1
*.iopin n8
*.iopin n9
xcdum top ndum unitcap
xc0 top n0 unitcap
xc1_1_ top n1 unitcap
xc1_0_ top n1 unitcap
xc2_3_ top n2 unitcap
xc2_2_ top n2 unitcap
xc2_1_ top n2 unitcap
xc2_0_ top n2 unitcap
xc3_7_ top n3 unitcap
xc3_6_ top n3 unitcap
xc3_5_ top n3 unitcap
xc3_4_ top n3 unitcap
xc3_3_ top n3 unitcap
xc3_2_ top n3 unitcap
xc3_1_ top n3 unitcap
xc3_0_ top n3 unitcap
xc4_15_ top n4 unitcap
xc4_14_ top n4 unitcap
xc4_13_ top n4 unitcap
xc4_12_ top n4 unitcap
xc4_11_ top n4 unitcap
xc4_10_ top n4 unitcap
xc4_9_ top n4 unitcap
xc4_8_ top n4 unitcap
xc4_7_ top n4 unitcap
xc4_6_ top n4 unitcap
xc4_5_ top n4 unitcap
xc4_4_ top n4 unitcap
xc4_3_ top n4 unitcap
xc4_2_ top n4 unitcap
xc4_1_ top n4 unitcap
xc4_0_ top n4 unitcap
xc5_31_ top n5 unitcap
xc5_30_ top n5 unitcap
xc5_29_ top n5 unitcap
xc5_28_ top n5 unitcap
xc5_27_ top n5 unitcap
xc5_26_ top n5 unitcap
xc5_25_ top n5 unitcap
xc5_24_ top n5 unitcap
xc5_23_ top n5 unitcap
xc5_22_ top n5 unitcap
xc5_21_ top n5 unitcap
xc5_20_ top n5 unitcap
xc5_19_ top n5 unitcap
xc5_18_ top n5 unitcap
xc5_17_ top n5 unitcap
xc5_16_ top n5 unitcap
xc5_15_ top n5 unitcap
xc5_14_ top n5 unitcap
xc5_13_ top n5 unitcap
xc5_12_ top n5 unitcap
xc5_11_ top n5 unitcap
xc5_10_ top n5 unitcap
xc5_9_ top n5 unitcap
xc5_8_ top n5 unitcap
xc5_7_ top n5 unitcap
xc5_6_ top n5 unitcap
xc5_5_ top n5 unitcap
xc5_4_ top n5 unitcap
xc5_3_ top n5 unitcap
xc5_2_ top n5 unitcap
xc5_1_ top n5 unitcap
xc5_0_ top n5 unitcap
xc6_63_ top n6 unitcap
xc6_62_ top n6 unitcap
xc6_61_ top n6 unitcap
xc6_60_ top n6 unitcap
xc6_59_ top n6 unitcap
xc6_58_ top n6 unitcap
xc6_57_ top n6 unitcap
xc6_56_ top n6 unitcap
xc6_55_ top n6 unitcap
xc6_54_ top n6 unitcap
xc6_53_ top n6 unitcap
xc6_52_ top n6 unitcap
xc6_51_ top n6 unitcap
xc6_50_ top n6 unitcap
xc6_49_ top n6 unitcap
xc6_48_ top n6 unitcap
xc6_47_ top n6 unitcap
xc6_46_ top n6 unitcap
xc6_45_ top n6 unitcap
xc6_44_ top n6 unitcap
xc6_43_ top n6 unitcap
xc6_42_ top n6 unitcap
xc6_41_ top n6 unitcap
xc6_40_ top n6 unitcap
xc6_39_ top n6 unitcap
xc6_38_ top n6 unitcap
xc6_37_ top n6 unitcap
xc6_36_ top n6 unitcap
xc6_35_ top n6 unitcap
xc6_34_ top n6 unitcap
xc6_33_ top n6 unitcap
xc6_32_ top n6 unitcap
xc6_31_ top n6 unitcap
xc6_30_ top n6 unitcap
xc6_29_ top n6 unitcap
xc6_28_ top n6 unitcap
xc6_27_ top n6 unitcap
xc6_26_ top n6 unitcap
xc6_25_ top n6 unitcap
xc6_24_ top n6 unitcap
xc6_23_ top n6 unitcap
xc6_22_ top n6 unitcap
xc6_21_ top n6 unitcap
xc6_20_ top n6 unitcap
xc6_19_ top n6 unitcap
xc6_18_ top n6 unitcap
xc6_17_ top n6 unitcap
xc6_16_ top n6 unitcap
xc6_15_ top n6 unitcap
xc6_14_ top n6 unitcap
xc6_13_ top n6 unitcap
xc6_12_ top n6 unitcap
xc6_11_ top n6 unitcap
xc6_10_ top n6 unitcap
xc6_9_ top n6 unitcap
xc6_8_ top n6 unitcap
xc6_7_ top n6 unitcap
xc6_6_ top n6 unitcap
xc6_5_ top n6 unitcap
xc6_4_ top n6 unitcap
xc6_3_ top n6 unitcap
xc6_2_ top n6 unitcap
xc6_1_ top n6 unitcap
xc6_0_ top n6 unitcap
xc7_127_ top n7 unitcap
xc7_126_ top n7 unitcap
xc7_125_ top n7 unitcap
xc7_124_ top n7 unitcap
xc7_123_ top n7 unitcap
xc7_122_ top n7 unitcap
xc7_121_ top n7 unitcap
xc7_120_ top n7 unitcap
xc7_119_ top n7 unitcap
xc7_118_ top n7 unitcap
xc7_117_ top n7 unitcap
xc7_116_ top n7 unitcap
xc7_115_ top n7 unitcap
xc7_114_ top n7 unitcap
xc7_113_ top n7 unitcap
xc7_112_ top n7 unitcap
xc7_111_ top n7 unitcap
xc7_110_ top n7 unitcap
xc7_109_ top n7 unitcap
xc7_108_ top n7 unitcap
xc7_107_ top n7 unitcap
xc7_106_ top n7 unitcap
xc7_105_ top n7 unitcap
xc7_104_ top n7 unitcap
xc7_103_ top n7 unitcap
xc7_102_ top n7 unitcap
xc7_101_ top n7 unitcap
xc7_100_ top n7 unitcap
xc7_99_ top n7 unitcap
xc7_98_ top n7 unitcap
xc7_97_ top n7 unitcap
xc7_96_ top n7 unitcap
xc7_95_ top n7 unitcap
xc7_94_ top n7 unitcap
xc7_93_ top n7 unitcap
xc7_92_ top n7 unitcap
xc7_91_ top n7 unitcap
xc7_90_ top n7 unitcap
xc7_89_ top n7 unitcap
xc7_88_ top n7 unitcap
xc7_87_ top n7 unitcap
xc7_86_ top n7 unitcap
xc7_85_ top n7 unitcap
xc7_84_ top n7 unitcap
xc7_83_ top n7 unitcap
xc7_82_ top n7 unitcap
xc7_81_ top n7 unitcap
xc7_80_ top n7 unitcap
xc7_79_ top n7 unitcap
xc7_78_ top n7 unitcap
xc7_77_ top n7 unitcap
xc7_76_ top n7 unitcap
xc7_75_ top n7 unitcap
xc7_74_ top n7 unitcap
xc7_73_ top n7 unitcap
xc7_72_ top n7 unitcap
xc7_71_ top n7 unitcap
xc7_70_ top n7 unitcap
xc7_69_ top n7 unitcap
xc7_68_ top n7 unitcap
xc7_67_ top n7 unitcap
xc7_66_ top n7 unitcap
xc7_65_ top n7 unitcap
xc7_64_ top n7 unitcap
xc7_63_ top n7 unitcap
xc7_62_ top n7 unitcap
xc7_61_ top n7 unitcap
xc7_60_ top n7 unitcap
xc7_59_ top n7 unitcap
xc7_58_ top n7 unitcap
xc7_57_ top n7 unitcap
xc7_56_ top n7 unitcap
xc7_55_ top n7 unitcap
xc7_54_ top n7 unitcap
xc7_53_ top n7 unitcap
xc7_52_ top n7 unitcap
xc7_51_ top n7 unitcap
xc7_50_ top n7 unitcap
xc7_49_ top n7 unitcap
xc7_48_ top n7 unitcap
xc7_47_ top n7 unitcap
xc7_46_ top n7 unitcap
xc7_45_ top n7 unitcap
xc7_44_ top n7 unitcap
xc7_43_ top n7 unitcap
xc7_42_ top n7 unitcap
xc7_41_ top n7 unitcap
xc7_40_ top n7 unitcap
xc7_39_ top n7 unitcap
xc7_38_ top n7 unitcap
xc7_37_ top n7 unitcap
xc7_36_ top n7 unitcap
xc7_35_ top n7 unitcap
xc7_34_ top n7 unitcap
xc7_33_ top n7 unitcap
xc7_32_ top n7 unitcap
xc7_31_ top n7 unitcap
xc7_30_ top n7 unitcap
xc7_29_ top n7 unitcap
xc7_28_ top n7 unitcap
xc7_27_ top n7 unitcap
xc7_26_ top n7 unitcap
xc7_25_ top n7 unitcap
xc7_24_ top n7 unitcap
xc7_23_ top n7 unitcap
xc7_22_ top n7 unitcap
xc7_21_ top n7 unitcap
xc7_20_ top n7 unitcap
xc7_19_ top n7 unitcap
xc7_18_ top n7 unitcap
xc7_17_ top n7 unitcap
xc7_16_ top n7 unitcap
xc7_15_ top n7 unitcap
xc7_14_ top n7 unitcap
xc7_13_ top n7 unitcap
xc7_12_ top n7 unitcap
xc7_11_ top n7 unitcap
xc7_10_ top n7 unitcap
xc7_9_ top n7 unitcap
xc7_8_ top n7 unitcap
xc7_7_ top n7 unitcap
xc7_6_ top n7 unitcap
xc7_5_ top n7 unitcap
xc7_4_ top n7 unitcap
xc7_3_ top n7 unitcap
xc7_2_ top n7 unitcap
xc7_1_ top n7 unitcap
xc7_0_ top n7 unitcap
xc8_255_ top n8 unitcap
xc8_254_ top n8 unitcap
xc8_253_ top n8 unitcap
xc8_252_ top n8 unitcap
xc8_251_ top n8 unitcap
xc8_250_ top n8 unitcap
xc8_249_ top n8 unitcap
xc8_248_ top n8 unitcap
xc8_247_ top n8 unitcap
xc8_246_ top n8 unitcap
xc8_245_ top n8 unitcap
xc8_244_ top n8 unitcap
xc8_243_ top n8 unitcap
xc8_242_ top n8 unitcap
xc8_241_ top n8 unitcap
xc8_240_ top n8 unitcap
xc8_239_ top n8 unitcap
xc8_238_ top n8 unitcap
xc8_237_ top n8 unitcap
xc8_236_ top n8 unitcap
xc8_235_ top n8 unitcap
xc8_234_ top n8 unitcap
xc8_233_ top n8 unitcap
xc8_232_ top n8 unitcap
xc8_231_ top n8 unitcap
xc8_230_ top n8 unitcap
xc8_229_ top n8 unitcap
xc8_228_ top n8 unitcap
xc8_227_ top n8 unitcap
xc8_226_ top n8 unitcap
xc8_225_ top n8 unitcap
xc8_224_ top n8 unitcap
xc8_223_ top n8 unitcap
xc8_222_ top n8 unitcap
xc8_221_ top n8 unitcap
xc8_220_ top n8 unitcap
xc8_219_ top n8 unitcap
xc8_218_ top n8 unitcap
xc8_217_ top n8 unitcap
xc8_216_ top n8 unitcap
xc8_215_ top n8 unitcap
xc8_214_ top n8 unitcap
xc8_213_ top n8 unitcap
xc8_212_ top n8 unitcap
xc8_211_ top n8 unitcap
xc8_210_ top n8 unitcap
xc8_209_ top n8 unitcap
xc8_208_ top n8 unitcap
xc8_207_ top n8 unitcap
xc8_206_ top n8 unitcap
xc8_205_ top n8 unitcap
xc8_204_ top n8 unitcap
xc8_203_ top n8 unitcap
xc8_202_ top n8 unitcap
xc8_201_ top n8 unitcap
xc8_200_ top n8 unitcap
xc8_199_ top n8 unitcap
xc8_198_ top n8 unitcap
xc8_197_ top n8 unitcap
xc8_196_ top n8 unitcap
xc8_195_ top n8 unitcap
xc8_194_ top n8 unitcap
xc8_193_ top n8 unitcap
xc8_192_ top n8 unitcap
xc8_191_ top n8 unitcap
xc8_190_ top n8 unitcap
xc8_189_ top n8 unitcap
xc8_188_ top n8 unitcap
xc8_187_ top n8 unitcap
xc8_186_ top n8 unitcap
xc8_185_ top n8 unitcap
xc8_184_ top n8 unitcap
xc8_183_ top n8 unitcap
xc8_182_ top n8 unitcap
xc8_181_ top n8 unitcap
xc8_180_ top n8 unitcap
xc8_179_ top n8 unitcap
xc8_178_ top n8 unitcap
xc8_177_ top n8 unitcap
xc8_176_ top n8 unitcap
xc8_175_ top n8 unitcap
xc8_174_ top n8 unitcap
xc8_173_ top n8 unitcap
xc8_172_ top n8 unitcap
xc8_171_ top n8 unitcap
xc8_170_ top n8 unitcap
xc8_169_ top n8 unitcap
xc8_168_ top n8 unitcap
xc8_167_ top n8 unitcap
xc8_166_ top n8 unitcap
xc8_165_ top n8 unitcap
xc8_164_ top n8 unitcap
xc8_163_ top n8 unitcap
xc8_162_ top n8 unitcap
xc8_161_ top n8 unitcap
xc8_160_ top n8 unitcap
xc8_159_ top n8 unitcap
xc8_158_ top n8 unitcap
xc8_157_ top n8 unitcap
xc8_156_ top n8 unitcap
xc8_155_ top n8 unitcap
xc8_154_ top n8 unitcap
xc8_153_ top n8 unitcap
xc8_152_ top n8 unitcap
xc8_151_ top n8 unitcap
xc8_150_ top n8 unitcap
xc8_149_ top n8 unitcap
xc8_148_ top n8 unitcap
xc8_147_ top n8 unitcap
xc8_146_ top n8 unitcap
xc8_145_ top n8 unitcap
xc8_144_ top n8 unitcap
xc8_143_ top n8 unitcap
xc8_142_ top n8 unitcap
xc8_141_ top n8 unitcap
xc8_140_ top n8 unitcap
xc8_139_ top n8 unitcap
xc8_138_ top n8 unitcap
xc8_137_ top n8 unitcap
xc8_136_ top n8 unitcap
xc8_135_ top n8 unitcap
xc8_134_ top n8 unitcap
xc8_133_ top n8 unitcap
xc8_132_ top n8 unitcap
xc8_131_ top n8 unitcap
xc8_130_ top n8 unitcap
xc8_129_ top n8 unitcap
xc8_128_ top n8 unitcap
xc8_127_ top n8 unitcap
xc8_126_ top n8 unitcap
xc8_125_ top n8 unitcap
xc8_124_ top n8 unitcap
xc8_123_ top n8 unitcap
xc8_122_ top n8 unitcap
xc8_121_ top n8 unitcap
xc8_120_ top n8 unitcap
xc8_119_ top n8 unitcap
xc8_118_ top n8 unitcap
xc8_117_ top n8 unitcap
xc8_116_ top n8 unitcap
xc8_115_ top n8 unitcap
xc8_114_ top n8 unitcap
xc8_113_ top n8 unitcap
xc8_112_ top n8 unitcap
xc8_111_ top n8 unitcap
xc8_110_ top n8 unitcap
xc8_109_ top n8 unitcap
xc8_108_ top n8 unitcap
xc8_107_ top n8 unitcap
xc8_106_ top n8 unitcap
xc8_105_ top n8 unitcap
xc8_104_ top n8 unitcap
xc8_103_ top n8 unitcap
xc8_102_ top n8 unitcap
xc8_101_ top n8 unitcap
xc8_100_ top n8 unitcap
xc8_99_ top n8 unitcap
xc8_98_ top n8 unitcap
xc8_97_ top n8 unitcap
xc8_96_ top n8 unitcap
xc8_95_ top n8 unitcap
xc8_94_ top n8 unitcap
xc8_93_ top n8 unitcap
xc8_92_ top n8 unitcap
xc8_91_ top n8 unitcap
xc8_90_ top n8 unitcap
xc8_89_ top n8 unitcap
xc8_88_ top n8 unitcap
xc8_87_ top n8 unitcap
xc8_86_ top n8 unitcap
xc8_85_ top n8 unitcap
xc8_84_ top n8 unitcap
xc8_83_ top n8 unitcap
xc8_82_ top n8 unitcap
xc8_81_ top n8 unitcap
xc8_80_ top n8 unitcap
xc8_79_ top n8 unitcap
xc8_78_ top n8 unitcap
xc8_77_ top n8 unitcap
xc8_76_ top n8 unitcap
xc8_75_ top n8 unitcap
xc8_74_ top n8 unitcap
xc8_73_ top n8 unitcap
xc8_72_ top n8 unitcap
xc8_71_ top n8 unitcap
xc8_70_ top n8 unitcap
xc8_69_ top n8 unitcap
xc8_68_ top n8 unitcap
xc8_67_ top n8 unitcap
xc8_66_ top n8 unitcap
xc8_65_ top n8 unitcap
xc8_64_ top n8 unitcap
xc8_63_ top n8 unitcap
xc8_62_ top n8 unitcap
xc8_61_ top n8 unitcap
xc8_60_ top n8 unitcap
xc8_59_ top n8 unitcap
xc8_58_ top n8 unitcap
xc8_57_ top n8 unitcap
xc8_56_ top n8 unitcap
xc8_55_ top n8 unitcap
xc8_54_ top n8 unitcap
xc8_53_ top n8 unitcap
xc8_52_ top n8 unitcap
xc8_51_ top n8 unitcap
xc8_50_ top n8 unitcap
xc8_49_ top n8 unitcap
xc8_48_ top n8 unitcap
xc8_47_ top n8 unitcap
xc8_46_ top n8 unitcap
xc8_45_ top n8 unitcap
xc8_44_ top n8 unitcap
xc8_43_ top n8 unitcap
xc8_42_ top n8 unitcap
xc8_41_ top n8 unitcap
xc8_40_ top n8 unitcap
xc8_39_ top n8 unitcap
xc8_38_ top n8 unitcap
xc8_37_ top n8 unitcap
xc8_36_ top n8 unitcap
xc8_35_ top n8 unitcap
xc8_34_ top n8 unitcap
xc8_33_ top n8 unitcap
xc8_32_ top n8 unitcap
xc8_31_ top n8 unitcap
xc8_30_ top n8 unitcap
xc8_29_ top n8 unitcap
xc8_28_ top n8 unitcap
xc8_27_ top n8 unitcap
xc8_26_ top n8 unitcap
xc8_25_ top n8 unitcap
xc8_24_ top n8 unitcap
xc8_23_ top n8 unitcap
xc8_22_ top n8 unitcap
xc8_21_ top n8 unitcap
xc8_20_ top n8 unitcap
xc8_19_ top n8 unitcap
xc8_18_ top n8 unitcap
xc8_17_ top n8 unitcap
xc8_16_ top n8 unitcap
xc8_15_ top n8 unitcap
xc8_14_ top n8 unitcap
xc8_13_ top n8 unitcap
xc8_12_ top n8 unitcap
xc8_11_ top n8 unitcap
xc8_10_ top n8 unitcap
xc8_9_ top n8 unitcap
xc8_8_ top n8 unitcap
xc8_7_ top n8 unitcap
xc8_6_ top n8 unitcap
xc8_5_ top n8 unitcap
xc8_4_ top n8 unitcap
xc8_3_ top n8 unitcap
xc8_2_ top n8 unitcap
xc8_1_ top n8 unitcap
xc8_0_ top n8 unitcap
xc9_511_ top n9 unitcap
xc9_510_ top n9 unitcap
xc9_509_ top n9 unitcap
xc9_508_ top n9 unitcap
xc9_507_ top n9 unitcap
xc9_506_ top n9 unitcap
xc9_505_ top n9 unitcap
xc9_504_ top n9 unitcap
xc9_503_ top n9 unitcap
xc9_502_ top n9 unitcap
xc9_501_ top n9 unitcap
xc9_500_ top n9 unitcap
xc9_499_ top n9 unitcap
xc9_498_ top n9 unitcap
xc9_497_ top n9 unitcap
xc9_496_ top n9 unitcap
xc9_495_ top n9 unitcap
xc9_494_ top n9 unitcap
xc9_493_ top n9 unitcap
xc9_492_ top n9 unitcap
xc9_491_ top n9 unitcap
xc9_490_ top n9 unitcap
xc9_489_ top n9 unitcap
xc9_488_ top n9 unitcap
xc9_487_ top n9 unitcap
xc9_486_ top n9 unitcap
xc9_485_ top n9 unitcap
xc9_484_ top n9 unitcap
xc9_483_ top n9 unitcap
xc9_482_ top n9 unitcap
xc9_481_ top n9 unitcap
xc9_480_ top n9 unitcap
xc9_479_ top n9 unitcap
xc9_478_ top n9 unitcap
xc9_477_ top n9 unitcap
xc9_476_ top n9 unitcap
xc9_475_ top n9 unitcap
xc9_474_ top n9 unitcap
xc9_473_ top n9 unitcap
xc9_472_ top n9 unitcap
xc9_471_ top n9 unitcap
xc9_470_ top n9 unitcap
xc9_469_ top n9 unitcap
xc9_468_ top n9 unitcap
xc9_467_ top n9 unitcap
xc9_466_ top n9 unitcap
xc9_465_ top n9 unitcap
xc9_464_ top n9 unitcap
xc9_463_ top n9 unitcap
xc9_462_ top n9 unitcap
xc9_461_ top n9 unitcap
xc9_460_ top n9 unitcap
xc9_459_ top n9 unitcap
xc9_458_ top n9 unitcap
xc9_457_ top n9 unitcap
xc9_456_ top n9 unitcap
xc9_455_ top n9 unitcap
xc9_454_ top n9 unitcap
xc9_453_ top n9 unitcap
xc9_452_ top n9 unitcap
xc9_451_ top n9 unitcap
xc9_450_ top n9 unitcap
xc9_449_ top n9 unitcap
xc9_448_ top n9 unitcap
xc9_447_ top n9 unitcap
xc9_446_ top n9 unitcap
xc9_445_ top n9 unitcap
xc9_444_ top n9 unitcap
xc9_443_ top n9 unitcap
xc9_442_ top n9 unitcap
xc9_441_ top n9 unitcap
xc9_440_ top n9 unitcap
xc9_439_ top n9 unitcap
xc9_438_ top n9 unitcap
xc9_437_ top n9 unitcap
xc9_436_ top n9 unitcap
xc9_435_ top n9 unitcap
xc9_434_ top n9 unitcap
xc9_433_ top n9 unitcap
xc9_432_ top n9 unitcap
xc9_431_ top n9 unitcap
xc9_430_ top n9 unitcap
xc9_429_ top n9 unitcap
xc9_428_ top n9 unitcap
xc9_427_ top n9 unitcap
xc9_426_ top n9 unitcap
xc9_425_ top n9 unitcap
xc9_424_ top n9 unitcap
xc9_423_ top n9 unitcap
xc9_422_ top n9 unitcap
xc9_421_ top n9 unitcap
xc9_420_ top n9 unitcap
xc9_419_ top n9 unitcap
xc9_418_ top n9 unitcap
xc9_417_ top n9 unitcap
xc9_416_ top n9 unitcap
xc9_415_ top n9 unitcap
xc9_414_ top n9 unitcap
xc9_413_ top n9 unitcap
xc9_412_ top n9 unitcap
xc9_411_ top n9 unitcap
xc9_410_ top n9 unitcap
xc9_409_ top n9 unitcap
xc9_408_ top n9 unitcap
xc9_407_ top n9 unitcap
xc9_406_ top n9 unitcap
xc9_405_ top n9 unitcap
xc9_404_ top n9 unitcap
xc9_403_ top n9 unitcap
xc9_402_ top n9 unitcap
xc9_401_ top n9 unitcap
xc9_400_ top n9 unitcap
xc9_399_ top n9 unitcap
xc9_398_ top n9 unitcap
xc9_397_ top n9 unitcap
xc9_396_ top n9 unitcap
xc9_395_ top n9 unitcap
xc9_394_ top n9 unitcap
xc9_393_ top n9 unitcap
xc9_392_ top n9 unitcap
xc9_391_ top n9 unitcap
xc9_390_ top n9 unitcap
xc9_389_ top n9 unitcap
xc9_388_ top n9 unitcap
xc9_387_ top n9 unitcap
xc9_386_ top n9 unitcap
xc9_385_ top n9 unitcap
xc9_384_ top n9 unitcap
xc9_383_ top n9 unitcap
xc9_382_ top n9 unitcap
xc9_381_ top n9 unitcap
xc9_380_ top n9 unitcap
xc9_379_ top n9 unitcap
xc9_378_ top n9 unitcap
xc9_377_ top n9 unitcap
xc9_376_ top n9 unitcap
xc9_375_ top n9 unitcap
xc9_374_ top n9 unitcap
xc9_373_ top n9 unitcap
xc9_372_ top n9 unitcap
xc9_371_ top n9 unitcap
xc9_370_ top n9 unitcap
xc9_369_ top n9 unitcap
xc9_368_ top n9 unitcap
xc9_367_ top n9 unitcap
xc9_366_ top n9 unitcap
xc9_365_ top n9 unitcap
xc9_364_ top n9 unitcap
xc9_363_ top n9 unitcap
xc9_362_ top n9 unitcap
xc9_361_ top n9 unitcap
xc9_360_ top n9 unitcap
xc9_359_ top n9 unitcap
xc9_358_ top n9 unitcap
xc9_357_ top n9 unitcap
xc9_356_ top n9 unitcap
xc9_355_ top n9 unitcap
xc9_354_ top n9 unitcap
xc9_353_ top n9 unitcap
xc9_352_ top n9 unitcap
xc9_351_ top n9 unitcap
xc9_350_ top n9 unitcap
xc9_349_ top n9 unitcap
xc9_348_ top n9 unitcap
xc9_347_ top n9 unitcap
xc9_346_ top n9 unitcap
xc9_345_ top n9 unitcap
xc9_344_ top n9 unitcap
xc9_343_ top n9 unitcap
xc9_342_ top n9 unitcap
xc9_341_ top n9 unitcap
xc9_340_ top n9 unitcap
xc9_339_ top n9 unitcap
xc9_338_ top n9 unitcap
xc9_337_ top n9 unitcap
xc9_336_ top n9 unitcap
xc9_335_ top n9 unitcap
xc9_334_ top n9 unitcap
xc9_333_ top n9 unitcap
xc9_332_ top n9 unitcap
xc9_331_ top n9 unitcap
xc9_330_ top n9 unitcap
xc9_329_ top n9 unitcap
xc9_328_ top n9 unitcap
xc9_327_ top n9 unitcap
xc9_326_ top n9 unitcap
xc9_325_ top n9 unitcap
xc9_324_ top n9 unitcap
xc9_323_ top n9 unitcap
xc9_322_ top n9 unitcap
xc9_321_ top n9 unitcap
xc9_320_ top n9 unitcap
xc9_319_ top n9 unitcap
xc9_318_ top n9 unitcap
xc9_317_ top n9 unitcap
xc9_316_ top n9 unitcap
xc9_315_ top n9 unitcap
xc9_314_ top n9 unitcap
xc9_313_ top n9 unitcap
xc9_312_ top n9 unitcap
xc9_311_ top n9 unitcap
xc9_310_ top n9 unitcap
xc9_309_ top n9 unitcap
xc9_308_ top n9 unitcap
xc9_307_ top n9 unitcap
xc9_306_ top n9 unitcap
xc9_305_ top n9 unitcap
xc9_304_ top n9 unitcap
xc9_303_ top n9 unitcap
xc9_302_ top n9 unitcap
xc9_301_ top n9 unitcap
xc9_300_ top n9 unitcap
xc9_299_ top n9 unitcap
xc9_298_ top n9 unitcap
xc9_297_ top n9 unitcap
xc9_296_ top n9 unitcap
xc9_295_ top n9 unitcap
xc9_294_ top n9 unitcap
xc9_293_ top n9 unitcap
xc9_292_ top n9 unitcap
xc9_291_ top n9 unitcap
xc9_290_ top n9 unitcap
xc9_289_ top n9 unitcap
xc9_288_ top n9 unitcap
xc9_287_ top n9 unitcap
xc9_286_ top n9 unitcap
xc9_285_ top n9 unitcap
xc9_284_ top n9 unitcap
xc9_283_ top n9 unitcap
xc9_282_ top n9 unitcap
xc9_281_ top n9 unitcap
xc9_280_ top n9 unitcap
xc9_279_ top n9 unitcap
xc9_278_ top n9 unitcap
xc9_277_ top n9 unitcap
xc9_276_ top n9 unitcap
xc9_275_ top n9 unitcap
xc9_274_ top n9 unitcap
xc9_273_ top n9 unitcap
xc9_272_ top n9 unitcap
xc9_271_ top n9 unitcap
xc9_270_ top n9 unitcap
xc9_269_ top n9 unitcap
xc9_268_ top n9 unitcap
xc9_267_ top n9 unitcap
xc9_266_ top n9 unitcap
xc9_265_ top n9 unitcap
xc9_264_ top n9 unitcap
xc9_263_ top n9 unitcap
xc9_262_ top n9 unitcap
xc9_261_ top n9 unitcap
xc9_260_ top n9 unitcap
xc9_259_ top n9 unitcap
xc9_258_ top n9 unitcap
xc9_257_ top n9 unitcap
xc9_256_ top n9 unitcap
xc9_255_ top n9 unitcap
xc9_254_ top n9 unitcap
xc9_253_ top n9 unitcap
xc9_252_ top n9 unitcap
xc9_251_ top n9 unitcap
xc9_250_ top n9 unitcap
xc9_249_ top n9 unitcap
xc9_248_ top n9 unitcap
xc9_247_ top n9 unitcap
xc9_246_ top n9 unitcap
xc9_245_ top n9 unitcap
xc9_244_ top n9 unitcap
xc9_243_ top n9 unitcap
xc9_242_ top n9 unitcap
xc9_241_ top n9 unitcap
xc9_240_ top n9 unitcap
xc9_239_ top n9 unitcap
xc9_238_ top n9 unitcap
xc9_237_ top n9 unitcap
xc9_236_ top n9 unitcap
xc9_235_ top n9 unitcap
xc9_234_ top n9 unitcap
xc9_233_ top n9 unitcap
xc9_232_ top n9 unitcap
xc9_231_ top n9 unitcap
xc9_230_ top n9 unitcap
xc9_229_ top n9 unitcap
xc9_228_ top n9 unitcap
xc9_227_ top n9 unitcap
xc9_226_ top n9 unitcap
xc9_225_ top n9 unitcap
xc9_224_ top n9 unitcap
xc9_223_ top n9 unitcap
xc9_222_ top n9 unitcap
xc9_221_ top n9 unitcap
xc9_220_ top n9 unitcap
xc9_219_ top n9 unitcap
xc9_218_ top n9 unitcap
xc9_217_ top n9 unitcap
xc9_216_ top n9 unitcap
xc9_215_ top n9 unitcap
xc9_214_ top n9 unitcap
xc9_213_ top n9 unitcap
xc9_212_ top n9 unitcap
xc9_211_ top n9 unitcap
xc9_210_ top n9 unitcap
xc9_209_ top n9 unitcap
xc9_208_ top n9 unitcap
xc9_207_ top n9 unitcap
xc9_206_ top n9 unitcap
xc9_205_ top n9 unitcap
xc9_204_ top n9 unitcap
xc9_203_ top n9 unitcap
xc9_202_ top n9 unitcap
xc9_201_ top n9 unitcap
xc9_200_ top n9 unitcap
xc9_199_ top n9 unitcap
xc9_198_ top n9 unitcap
xc9_197_ top n9 unitcap
xc9_196_ top n9 unitcap
xc9_195_ top n9 unitcap
xc9_194_ top n9 unitcap
xc9_193_ top n9 unitcap
xc9_192_ top n9 unitcap
xc9_191_ top n9 unitcap
xc9_190_ top n9 unitcap
xc9_189_ top n9 unitcap
xc9_188_ top n9 unitcap
xc9_187_ top n9 unitcap
xc9_186_ top n9 unitcap
xc9_185_ top n9 unitcap
xc9_184_ top n9 unitcap
xc9_183_ top n9 unitcap
xc9_182_ top n9 unitcap
xc9_181_ top n9 unitcap
xc9_180_ top n9 unitcap
xc9_179_ top n9 unitcap
xc9_178_ top n9 unitcap
xc9_177_ top n9 unitcap
xc9_176_ top n9 unitcap
xc9_175_ top n9 unitcap
xc9_174_ top n9 unitcap
xc9_173_ top n9 unitcap
xc9_172_ top n9 unitcap
xc9_171_ top n9 unitcap
xc9_170_ top n9 unitcap
xc9_169_ top n9 unitcap
xc9_168_ top n9 unitcap
xc9_167_ top n9 unitcap
xc9_166_ top n9 unitcap
xc9_165_ top n9 unitcap
xc9_164_ top n9 unitcap
xc9_163_ top n9 unitcap
xc9_162_ top n9 unitcap
xc9_161_ top n9 unitcap
xc9_160_ top n9 unitcap
xc9_159_ top n9 unitcap
xc9_158_ top n9 unitcap
xc9_157_ top n9 unitcap
xc9_156_ top n9 unitcap
xc9_155_ top n9 unitcap
xc9_154_ top n9 unitcap
xc9_153_ top n9 unitcap
xc9_152_ top n9 unitcap
xc9_151_ top n9 unitcap
xc9_150_ top n9 unitcap
xc9_149_ top n9 unitcap
xc9_148_ top n9 unitcap
xc9_147_ top n9 unitcap
xc9_146_ top n9 unitcap
xc9_145_ top n9 unitcap
xc9_144_ top n9 unitcap
xc9_143_ top n9 unitcap
xc9_142_ top n9 unitcap
xc9_141_ top n9 unitcap
xc9_140_ top n9 unitcap
xc9_139_ top n9 unitcap
xc9_138_ top n9 unitcap
xc9_137_ top n9 unitcap
xc9_136_ top n9 unitcap
xc9_135_ top n9 unitcap
xc9_134_ top n9 unitcap
xc9_133_ top n9 unitcap
xc9_132_ top n9 unitcap
xc9_131_ top n9 unitcap
xc9_130_ top n9 unitcap
xc9_129_ top n9 unitcap
xc9_128_ top n9 unitcap
xc9_127_ top n9 unitcap
xc9_126_ top n9 unitcap
xc9_125_ top n9 unitcap
xc9_124_ top n9 unitcap
xc9_123_ top n9 unitcap
xc9_122_ top n9 unitcap
xc9_121_ top n9 unitcap
xc9_120_ top n9 unitcap
xc9_119_ top n9 unitcap
xc9_118_ top n9 unitcap
xc9_117_ top n9 unitcap
xc9_116_ top n9 unitcap
xc9_115_ top n9 unitcap
xc9_114_ top n9 unitcap
xc9_113_ top n9 unitcap
xc9_112_ top n9 unitcap
xc9_111_ top n9 unitcap
xc9_110_ top n9 unitcap
xc9_109_ top n9 unitcap
xc9_108_ top n9 unitcap
xc9_107_ top n9 unitcap
xc9_106_ top n9 unitcap
xc9_105_ top n9 unitcap
xc9_104_ top n9 unitcap
xc9_103_ top n9 unitcap
xc9_102_ top n9 unitcap
xc9_101_ top n9 unitcap
xc9_100_ top n9 unitcap
xc9_99_ top n9 unitcap
xc9_98_ top n9 unitcap
xc9_97_ top n9 unitcap
xc9_96_ top n9 unitcap
xc9_95_ top n9 unitcap
xc9_94_ top n9 unitcap
xc9_93_ top n9 unitcap
xc9_92_ top n9 unitcap
xc9_91_ top n9 unitcap
xc9_90_ top n9 unitcap
xc9_89_ top n9 unitcap
xc9_88_ top n9 unitcap
xc9_87_ top n9 unitcap
xc9_86_ top n9 unitcap
xc9_85_ top n9 unitcap
xc9_84_ top n9 unitcap
xc9_83_ top n9 unitcap
xc9_82_ top n9 unitcap
xc9_81_ top n9 unitcap
xc9_80_ top n9 unitcap
xc9_79_ top n9 unitcap
xc9_78_ top n9 unitcap
xc9_77_ top n9 unitcap
xc9_76_ top n9 unitcap
xc9_75_ top n9 unitcap
xc9_74_ top n9 unitcap
xc9_73_ top n9 unitcap
xc9_72_ top n9 unitcap
xc9_71_ top n9 unitcap
xc9_70_ top n9 unitcap
xc9_69_ top n9 unitcap
xc9_68_ top n9 unitcap
xc9_67_ top n9 unitcap
xc9_66_ top n9 unitcap
xc9_65_ top n9 unitcap
xc9_64_ top n9 unitcap
xc9_63_ top n9 unitcap
xc9_62_ top n9 unitcap
xc9_61_ top n9 unitcap
xc9_60_ top n9 unitcap
xc9_59_ top n9 unitcap
xc9_58_ top n9 unitcap
xc9_57_ top n9 unitcap
xc9_56_ top n9 unitcap
xc9_55_ top n9 unitcap
xc9_54_ top n9 unitcap
xc9_53_ top n9 unitcap
xc9_52_ top n9 unitcap
xc9_51_ top n9 unitcap
xc9_50_ top n9 unitcap
xc9_49_ top n9 unitcap
xc9_48_ top n9 unitcap
xc9_47_ top n9 unitcap
xc9_46_ top n9 unitcap
xc9_45_ top n9 unitcap
xc9_44_ top n9 unitcap
xc9_43_ top n9 unitcap
xc9_42_ top n9 unitcap
xc9_41_ top n9 unitcap
xc9_40_ top n9 unitcap
xc9_39_ top n9 unitcap
xc9_38_ top n9 unitcap
xc9_37_ top n9 unitcap
xc9_36_ top n9 unitcap
xc9_35_ top n9 unitcap
xc9_34_ top n9 unitcap
xc9_33_ top n9 unitcap
xc9_32_ top n9 unitcap
xc9_31_ top n9 unitcap
xc9_30_ top n9 unitcap
xc9_29_ top n9 unitcap
xc9_28_ top n9 unitcap
xc9_27_ top n9 unitcap
xc9_26_ top n9 unitcap
xc9_25_ top n9 unitcap
xc9_24_ top n9 unitcap
xc9_23_ top n9 unitcap
xc9_22_ top n9 unitcap
xc9_21_ top n9 unitcap
xc9_20_ top n9 unitcap
xc9_19_ top n9 unitcap
xc9_18_ top n9 unitcap
xc9_17_ top n9 unitcap
xc9_16_ top n9 unitcap
xc9_15_ top n9 unitcap
xc9_14_ top n9 unitcap
xc9_13_ top n9 unitcap
xc9_12_ top n9 unitcap
xc9_11_ top n9 unitcap
xc9_10_ top n9 unitcap
xc9_9_ top n9 unitcap
xc9_8_ top n9 unitcap
xc9_7_ top n9 unitcap
xc9_6_ top n9 unitcap
xc9_5_ top n9 unitcap
xc9_4_ top n9 unitcap
xc9_3_ top n9 unitcap
xc9_2_ top n9 unitcap
xc9_1_ top n9 unitcap
xc9_0_ top n9 unitcap
xegdedum_7_ top top unitcap
xegdedum_6_ top top unitcap
xegdedum_5_ top top unitcap
xegdedum_4_ top top unitcap
xegdedum_3_ top top unitcap
xegdedum_2_ top top unitcap
xegdedum_1_ top top unitcap
xegdedum_0_ top top unitcap
.ends


* expanding   symbol:  switches/bootstrapped_sw_hv.sym # of pins=5
* sym_path: /home/christoph/Studium/projekte/design/design/switches/bootstrapped_sw_hv.sym
* sch_path: /home/christoph/Studium/projekte/design/design/switches/bootstrapped_sw_hv.sch
.subckt bootstrapped_sw_hv  out en vdd in vss
*.iopin out
*.ipin en
*.iopin vss
*.iopin vdd
*.iopin in
xinv1 vdd en enb vss inv_lvt
XCbs_4_ vbsh vbsl sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XCbs_3_ vbsh vbsl sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XCbs_2_ vbsh vbsl sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XCbs_1_ vbsh vbsl sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XCbs_0_ vbsh vbsl sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XM3 vdd vg vbsh vbsh sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 vg enb vbsh vbsh sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMs out vg in vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 vbsl vg in vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 vbsl enb vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMs2 vss enb vs vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMs1 vs vdd vg vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  sar_10b/comparator/trim.sym # of pins=3
* sym_path: /home/christoph/Studium/projekte/design/design/sar_10b/comparator/trim.sym
* sch_path: /home/christoph/Studium/projekte/design/design/sar_10b/comparator/trim.sch
.subckt trim  drain d_4_ d_3_ d_2_ d_1_ d_0_ vss
*.iopin vss
*.ipin d_4_,d_3_,d_2_,d_1_,d_0_
*.opin drain
XM4_7_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4_6_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4_5_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4_4_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4_3_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4_2_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4_1_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4_0_ n4 d_4_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3_3_ n3 d_3_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3_2_ n3 d_3_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3_1_ n3 d_3_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3_0_ n3 d_3_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2_1_ n2 d_2_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2_0_ n2 d_2_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 n1 d_1_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM0 n0 d_0_ vss vss sky130_fd_pr__nfet_01v8_lvt L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
x4_7_ drain n4 trimcap
x4_6_ drain n4 trimcap
x4_5_ drain n4 trimcap
x4_4_ drain n4 trimcap
x4_3_ drain n4 trimcap
x4_2_ drain n4 trimcap
x4_1_ drain n4 trimcap
x4_0_ drain n4 trimcap
x3_3_ drain n3 trimcap
x3_2_ drain n3 trimcap
x3_1_ drain n3 trimcap
x3_0_ drain n3 trimcap
x2_1_ drain n2 trimcap
x2_0_ drain n2 trimcap
x1 drain n1 trimcap
x0 drain n0 trimcap
Cpar10 n1 n0 30e-18 m=1
Cpar43 n4 n3 30e-18 m=8
Cpar42 n4 n2 30e-18 m=4
Cpar41 n4 n1 30e-18 m=1
Cpar40 n4 n0 30e-18 m=1
.ends


* expanding   symbol:  bandgap/bg_res.sym # of pins=5
* sym_path: /home/christoph/Studium/projekte/design/design/bandgap/bg_res.sym
* sch_path: /home/christoph/Studium/projekte/design/design/bandgap/bg_res.sch
.subckt bg_res  b a d c vss
*.ipin a
*.ipin b
*.opin c
*.opin d
*.iopin vss
XR1 net1 a vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR2 net2 b vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR3 net6 net1 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR4 net5 net2 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR5 net3 net6 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR6 net4 net5 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR7 net10 net3 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR8 net9 net4 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR9 net7 net10 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR10 net8 net9 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR11 net12 net7 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR12 net11 net8 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR13 net14 net12 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR14 net13 net11 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR15 net16 net14 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR16 net15 net13 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR17 net18 net16 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR18 net17 net15 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR19 c net18 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
XR20 d net17 vss sky130_fd_pr__res_xhigh_po W=0.69 L=13 mult=1 m=1
.ends


* expanding   symbol:  bandgap/bg_trim.sym # of pins=4
* sym_path: /home/christoph/Studium/projekte/design/design/bandgap/bg_trim.sym
* sch_path: /home/christoph/Studium/projekte/design/design/bandgap/bg_trim.sch
.subckt bg_trim  top bot ctl_15_ ctl_14_ ctl_13_ ctl_12_ ctl_11_ ctl_10_ ctl_9_ ctl_8_ ctl_7_ ctl_6_
+ ctl_5_ ctl_4_ ctl_3_ ctl_2_ ctl_1_ ctl_0_ vss
*.iopin vss
*.ipin
*+ ctl_15_,ctl_14_,ctl_13_,ctl_12_,ctl_11_,ctl_10_,ctl_9_,ctl_8_,ctl_7_,ctl_6_,ctl_5_,ctl_4_,ctl_3_,ctl_2_,ctl_1_,ctl_0_
*.iopin bot
*.iopin top
XM0 net1 ctl_0_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM1 net2 ctl_1_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM2 net3 ctl_2_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM3 net4 ctl_3_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM4 net5 ctl_4_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM5 net6 ctl_5_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM6 net7 ctl_6_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM7 net8 ctl_7_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM12 net10 ctl_12_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM13 net11 ctl_13_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM14 net12 ctl_14_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM15 top ctl_15_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM8 net13 ctl_8_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM9 net14 ctl_9_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM10 net15 ctl_10_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XM11 net9 ctl_11_ bot vss sky130_fd_pr__nfet_01v8 L=0.5 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XR15 net12 top vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR1 net1 net2 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR2 net2 net3 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR3 net3 net4 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR4 net4 net5 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR5 net5 net6 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR6 net6 net7 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR7 net7 net8 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR8 net8 net13 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR9 net13 net14 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR10 net14 net15 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR11 net15 net9 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR12 net9 net10 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR13 net10 net11 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR14 net11 net12 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
XR16 bot net1 vss sky130_fd_pr__res_high_po W=1.41 L=2.8 mult=1 m=1
.ends


* expanding   symbol:  opamp/se_folded_cascode_p.sym # of pins=6
* sym_path: /home/christoph/Studium/projekte/design/design/opamp/se_folded_cascode_p.sym
* sch_path: /home/christoph/Studium/projekte/design/design/opamp/se_folded_cascode_p.sch
.subckt se_folded_cascode_p  vdd out inp inn vss bias
*.ipin inn
*.ipin inp
*.opin out
*.iopin bias
*.iopin vdd
*.iopin vss
XM3 out1p inn diff vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM2 out1n inp diff vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM1 diff vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM4 out1n vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM5 out1p vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM6 mirr vbn2 out1n vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM7 out vbn2 out1p vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM8 mirr bias nd10 vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM9 out bias nd11 vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM10 nd10 mirr vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM11 nd11 mirr vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XMB1 bias bias vbp1 vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XMB2 vbp1 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XMB3 vbn2 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XMB4 vbn2 vbn2 vbn1 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XMB5 vbn1 vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XMDUM1_41_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_40_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_39_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_38_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_37_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_36_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_35_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_34_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_33_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_32_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_31_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_30_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_29_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_28_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_27_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_26_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_25_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_24_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_23_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_22_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_21_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_20_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_19_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_18_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_17_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_16_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_15_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_14_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_13_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_12_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_11_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_10_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_9_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_8_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_7_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_6_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_5_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_4_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_3_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_2_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_1_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_0_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_3_ mirr mirr mirr vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_2_ mirr mirr mirr vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_1_ mirr mirr mirr vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_0_ mirr mirr mirr vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_3_ bias bias bias vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_2_ bias bias bias vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_1_ bias bias bias vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_0_ bias bias bias vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_23_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_22_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_21_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_20_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_19_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_18_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_17_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_16_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_15_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_14_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_13_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_12_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_11_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_10_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_9_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_8_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_7_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_6_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_5_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_4_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_3_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_2_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_1_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_0_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM5_3_ vbn2 vbn2 vbn2 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM5_2_ vbn2 vbn2 vbn2 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM5_1_ vbn2 vbn2 vbn2 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM5_0_ vbn2 vbn2 vbn2 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_43_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_42_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_41_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_40_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_39_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_38_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_37_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_36_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_35_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_34_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_33_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_32_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_31_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_30_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_29_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_28_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_27_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_26_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_25_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_24_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_23_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_22_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_21_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_20_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_19_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_18_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_17_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_16_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_15_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_14_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_13_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_12_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_11_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_10_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_9_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_8_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_7_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_6_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_5_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_4_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_3_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_2_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_1_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_0_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM7_3_ diff diff diff vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM7_2_ diff diff diff vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM7_1_ diff diff diff vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM7_0_ diff diff diff vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  bias/bias_amp.sym # of pins=6
* sym_path: /home/christoph/Studium/projekte/design/design/bias/bias_amp.sym
* sch_path: /home/christoph/Studium/projekte/design/design/bias/bias_amp.sch
.subckt bias_amp  vdd out inp inn vss bias
*.iopin vdd
*.iopin bias
*.ipin inp
*.ipin inn
*.opin out
*.iopin vss
XM3 mirr mirr vdd vdd sky130_fd_pr__pfet_01v8_lvt L=10 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM4 out mirr vdd vdd sky130_fd_pr__pfet_01v8_lvt L=10 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM1 mirr inp diff vss sky130_fd_pr__nfet_01v8_lvt L=8 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM2 out inn diff vss sky130_fd_pr__nfet_01v8_lvt L=8 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM5 net1 bias vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM6 bias bias vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XM5s diff bias net1 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
.ends


* expanding   symbol:  clkdiv/clkdiv.sym # of pins=5
* sym_path: /home/christoph/Studium/projekte/design/design/clkdiv/clkdiv.sym
* sch_path: /home/christoph/Studium/projekte/design/design/clkdiv/clkdiv.sch
.subckt clkdiv  dvss in out rst_b dvdd
*.ipin in
*.ipin rst_b
*.opin out
*.iopin dvdd
*.iopin dvss
x6 in net1 rst_b dvss dvss dvdd dvdd div2 net5 sky130_fd_sc_hd__dfrbp_1
x8 div2 dvss dvss dvdd dvdd net1 sky130_fd_sc_hd__inv_1
x1 div2 net2 rst_b dvss dvss dvdd dvdd div4 net6 sky130_fd_sc_hd__dfrbp_1
x2 div4 dvss dvss dvdd dvdd net2 sky130_fd_sc_hd__inv_1
x3 div4 net3 rst_b dvss dvss dvdd dvdd div8 net7 sky130_fd_sc_hd__dfrbp_1
x4 div8 dvss dvss dvdd dvdd net3 sky130_fd_sc_hd__inv_1
x5 div8 net4 rst_b dvss dvss dvdd dvdd out net8 sky130_fd_sc_hd__dfrbp_1
x7 out dvss dvss dvdd dvdd net4 sky130_fd_sc_hd__inv_1
xdec_7_ dvss dvss dvdd dvdd sky130_fd_sc_hd__decap_4
xdec_6_ dvss dvss dvdd dvdd sky130_fd_sc_hd__decap_4
xdec_5_ dvss dvss dvdd dvdd sky130_fd_sc_hd__decap_4
xdec_4_ dvss dvss dvdd dvdd sky130_fd_sc_hd__decap_4
xdec_3_ dvss dvss dvdd dvdd sky130_fd_sc_hd__decap_4
xdec_2_ dvss dvss dvdd dvdd sky130_fd_sc_hd__decap_4
xdec_1_ dvss dvss dvdd dvdd sky130_fd_sc_hd__decap_4
xdec_0_ dvss dvss dvdd dvdd sky130_fd_sc_hd__decap_4
xtap dvss dvdd sky130_fd_sc_hd__tapvpwrvgnd_1
.ends


* expanding   symbol:  switches/passgate.sym # of pins=5
* sym_path: /home/christoph/Studium/projekte/design/design/switches/passgate.sym
* sch_path: /home/christoph/Studium/projekte/design/design/switches/passgate.sch
.subckt passgate  out en vdd in vss
*.iopin out
*.ipin en
*.iopin vss
*.iopin vdd
*.iopin in
x2 vdd en enb vss inv_lvt
x1 vdd enb en_buf vss inv_lvt
XMSN out en_buf in vss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMSP in enb out vdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  testbuffer/mux.sym # of pins=5
* sym_path: /home/christoph/Studium/projekte/design/design/testbuffer/mux.sym
* sch_path: /home/christoph/Studium/projekte/design/design/testbuffer/mux.sch
.subckt mux  out vdd vss inp_7_ inp_6_ inp_5_ inp_4_ inp_3_ inp_2_ inp_1_ inp_0_ sel_2_ sel_1_
+ sel_0_
*.iopin out
*.ipin inp_7_,inp_6_,inp_5_,inp_4_,inp_3_,inp_2_,inp_1_,inp_0_
*.iopin vss
*.iopin vdd
*.ipin sel_2_,sel_1_,sel_0_
xpg1 out enm_1_ vdd inp_1_ vss passgate
xpg0 out enm_0_ vdd inp_0_ vss passgate
xpg3 out enm_3_ vdd inp_3_ vss passgate
xpg2 out enm_2_ vdd inp_2_ vss passgate
xpg5 out enm_5_ vdd inp_5_ vss passgate
xpg4 out enm_4_ vdd inp_4_ vss passgate
xpg6 out enm_6_ vdd inp_6_ vss passgate
xpg7 out enm_7_ vdd inp_7_ vss passgate
xdec enm_5_ vdd vss enm_4_ enm_3_ enm_2_ enm_1_ enm_0_ enm_6_ enm_7_ sel_0_ sel_1_ sel_2_
+ decoder3to8
.ends


* expanding   symbol:  opamp/se_folded_cascode_np_ab.sym # of pins=6
* sym_path: /home/christoph/Studium/projekte/design/design/opamp/se_folded_cascode_np_ab.sym
* sch_path: /home/christoph/Studium/projekte/design/design/opamp/se_folded_cascode_np_ab.sch
.subckt se_folded_cascode_np_ab  vdd out inp inn vss bias
*.iopin vdd
*.iopin bias
*.ipin inp
*.ipin inn
*.iopin vss
*.opin out
XM4 outa1n outa1n vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=12 m=12 
XM5 outa1p outa1n vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=12 m=12 
XMIN1 diffa vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=8 m=8 
XMB2 vbn1 vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XMB1 bias bias vbn1 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XMIN2 outa1n inn diffa vss sky130_fd_pr__nfet_01v8_lvt L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8 
XMIN3 outa1p inp diffa vss sky130_fd_pr__nfet_01v8_lvt L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8 
XMB5 vbp1 vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XM7 outs1 mirr outa1p vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM6 mirr mirr outa1n vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM8 mirr bias outb1n vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM9 outs1 bias outb1p vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XM10 outb1n vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=24 m=24 
XM11 outb1p vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=24 m=24 
XMB3 vbp2 vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XMB4 vbp2 vbp2 vbp1 vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XMIP2 outb1n inn diffb vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8 
XMIP3 outb1p inp diffb vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8 
XMIP1 diffb vbp1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=16 m=16 
XMON out outs1 vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XMOP out outs1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=4 m=4 
XC1_1_ out outs1 sky130_fd_pr__cap_mim_m3_1 W=25 L=25 MF=1 m=1
XC1_0_ out outs1 sky130_fd_pr__cap_mim_m3_1 W=25 L=25 MF=1 m=1
XMDUM6_3_ outs1 outs1 outs1 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_2_ outs1 outs1 outs1 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_1_ outs1 outs1 outs1 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM6_0_ outs1 outs1 outs1 vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM7_3_ mirr mirr mirr vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM7_2_ mirr mirr mirr vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM7_1_ mirr mirr mirr vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM7_0_ mirr mirr mirr vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_19_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_18_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_17_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_16_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_15_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_14_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_13_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_12_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_11_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_10_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_9_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_8_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_7_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_6_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_5_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_4_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_3_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_2_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_1_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM8_0_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=4 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_79_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_78_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_77_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_76_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_75_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_74_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_73_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_72_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_71_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_70_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_69_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_68_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_67_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_66_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_65_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_64_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_63_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_62_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_61_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_60_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_59_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_58_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_57_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_56_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_55_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_54_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_53_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_52_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_51_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_50_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_49_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_48_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_47_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_46_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_45_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_44_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_43_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_42_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_41_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_40_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_39_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_38_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_37_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_36_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_35_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_34_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_33_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_32_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_31_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_30_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_29_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_28_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_27_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_26_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_25_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_24_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_23_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_22_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_21_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_20_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_19_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_18_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_17_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_16_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_15_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_14_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_13_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_12_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_11_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_10_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_9_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_8_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_7_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_6_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_5_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_4_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_3_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_2_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_1_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM3_0_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_3_ mirr mirr mirr vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_2_ mirr mirr mirr vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_1_ mirr mirr mirr vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM4_0_ mirr mirr mirr vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM5_3_ outs1 outs1 outs1 vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM5_2_ outs1 outs1 outs1 vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM5_1_ outs1 outs1 outs1 vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM5_0_ outs1 outs1 outs1 vdd sky130_fd_pr__pfet_01v8_lvt L=4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM11 diffa diffa diffa vss sky130_fd_pr__nfet_01v8_lvt L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4 
XMDUM12 diffb diffb diffb vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4 
XMDUM9_35_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_34_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_33_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_32_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_31_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_30_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_29_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_28_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_27_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_26_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_25_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_24_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_23_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_22_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_21_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_20_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_19_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_18_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_17_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_16_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_15_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_14_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_13_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_12_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_11_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_10_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_9_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_8_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_7_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_6_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_5_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_4_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_3_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_2_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_1_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM9_0_ vss vss vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM10_7_ vss vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM10_6_ vss vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM10_5_ vss vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM10_4_ vss vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM10_3_ vss vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM10_2_ vss vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM10_1_ vss vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM10_0_ vss vbn1 vss vss sky130_fd_pr__nfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_27_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_26_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_25_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_24_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_23_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_22_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_21_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_20_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_19_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_18_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_17_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_16_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_15_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_14_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_13_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_12_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_11_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_10_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_9_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_8_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_7_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_6_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_5_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_4_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_3_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_2_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_1_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM1_0_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_31_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_30_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_29_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_28_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_27_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_26_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_25_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_24_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_23_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_22_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_21_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_20_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_19_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_18_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_17_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_16_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_15_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_14_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_13_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_12_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_11_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_10_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_9_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_8_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_7_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_6_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_5_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_4_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_3_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_2_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_1_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
XMDUM2_0_ vdd vdd vdd vdd sky130_fd_pr__pfet_01v8_lvt L=1 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 
.ends


* expanding   symbol:  sar_10b/unitcap/unitcap.sym # of pins=2
* sym_path: /home/christoph/Studium/projekte/design/design/sar_10b/unitcap/unitcap.sym
* sch_path: /home/christoph/Studium/projekte/design/design/sar_10b/unitcap/unitcap.sch
.subckt unitcap  cp cn
*.iopin cp
*.iopin cn
C1 cp cn 2.9f m=1
.ends


* expanding   symbol:  sar_10b/comparator/trimcap.sym # of pins=2
* sym_path: /home/christoph/Studium/projekte/design/design/sar_10b/comparator/trimcap.sym
* sch_path: /home/christoph/Studium/projekte/design/design/sar_10b/comparator/trimcap.sch
.subckt trimcap  cp cn
*.iopin cp
*.iopin cn
c0 cp cn 1.25f m=1
.ends
